* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
X_3155_ net541 net496 _2596_ VPWR VGND sg13g2_and2_1
XFILLER_39_299 VPWR VGND sg13g2_fill_1
X_3086_ VPWR _2527_ net522 VGND sg13g2_inv_1
XFILLER_35_450 VPWR VGND sg13g2_fill_1
XFILLER_36_951 VPWR VGND sg13g2_decap_8
X_3988_ _0959_ VPWR _0963_ VGND _0945_ _0960_ sg13g2_o21ai_1
XFILLER_11_829 VPWR VGND sg13g2_fill_1
X_5727_ net716 _2490_ net615 _2492_ VPWR VGND sg13g2_nand3_1
X_5658_ _2445_ mydesign.accum\[6\] _2446_ VPWR VGND sg13g2_xor2_1
X_5589_ _2381_ _2374_ _2380_ VPWR VGND sg13g2_nand2_1
X_4609_ net550 mydesign.inputs\[2\]\[16\] _1515_ VPWR VGND sg13g2_nor2_1
Xhold351 mydesign.accum\[11\] VPWR VGND net970 sg13g2_dlygate4sd3_1
Xhold362 mydesign.pe_inputs\[42\] VPWR VGND net981 sg13g2_dlygate4sd3_1
Xhold340 mydesign.accum\[58\] VPWR VGND net959 sg13g2_dlygate4sd3_1
Xhold384 mydesign.accum\[88\] VPWR VGND net1003 sg13g2_dlygate4sd3_1
X_5993__138 VPWR VGND net138 sg13g2_tiehi
Xhold395 _0232_ VPWR VGND net1014 sg13g2_dlygate4sd3_1
Xhold373 mydesign.accum\[19\] VPWR VGND net992 sg13g2_dlygate4sd3_1
XFILLER_46_726 VPWR VGND sg13g2_decap_8
XFILLER_45_247 VPWR VGND sg13g2_fill_1
XFILLER_26_41 VPWR VGND sg13g2_fill_2
XFILLER_27_962 VPWR VGND sg13g2_decap_8
XFILLER_42_954 VPWR VGND sg13g2_decap_8
XFILLER_14_645 VPWR VGND sg13g2_decap_4
XFILLER_41_486 VPWR VGND sg13g2_fill_1
XFILLER_10_840 VPWR VGND sg13g2_decap_8
XFILLER_6_822 VPWR VGND sg13g2_fill_2
X_5913__331 VPWR VGND net331 sg13g2_tiehi
X_4960_ _1815_ mydesign.pe_weights\[37\] mydesign.pe_inputs\[26\] VPWR VGND sg13g2_nand2_1
XFILLER_18_995 VPWR VGND sg13g2_decap_8
XFILLER_33_910 VPWR VGND sg13g2_decap_8
X_4891_ _1764_ net697 _1762_ VPWR VGND sg13g2_nand2_1
X_3911_ _0897_ _0883_ _0899_ VPWR VGND sg13g2_xor2_1
X_3842_ VGND VPWR net572 _0832_ _0126_ _0833_ sg13g2_a21oi_1
XFILLER_20_604 VPWR VGND sg13g2_fill_2
XFILLER_33_987 VPWR VGND sg13g2_decap_8
X_3773_ net622 VPWR _0775_ VGND net1076 net433 sg13g2_o21ai_1
X_5512_ _2314_ _2313_ _2312_ VPWR VGND sg13g2_nand2b_1
X_5443_ net477 VPWR _2249_ VGND net729 _2248_ sg13g2_o21ai_1
X_5374_ _2188_ mydesign.pe_inputs\[15\] mydesign.pe_weights\[25\] VPWR VGND sg13g2_nand2_1
X_4325_ net479 VPWR _1266_ VGND net580 net951 sg13g2_o21ai_1
X_4256_ _1198_ _1195_ _1200_ VPWR VGND sg13g2_xor2_1
X_4187_ _1144_ _1143_ _1141_ VPWR VGND sg13g2_nand2b_1
X_3207_ _2636_ VPWR _0011_ VGND _2518_ _2633_ sg13g2_o21ai_1
XFILLER_28_715 VPWR VGND sg13g2_fill_2
X_3138_ VPWR _2579_ net757 VGND sg13g2_inv_1
XFILLER_43_718 VPWR VGND sg13g2_decap_8
XFILLER_28_759 VPWR VGND sg13g2_fill_1
XFILLER_10_147 VPWR VGND sg13g2_fill_1
Xhold170 mydesign.pe_weights\[43\] VPWR VGND net789 sg13g2_dlygate4sd3_1
Xhold181 mydesign.inputs\[1\]\[11\] VPWR VGND net800 sg13g2_dlygate4sd3_1
Xhold192 mydesign.pe_weights\[45\] VPWR VGND net811 sg13g2_dlygate4sd3_1
XFILLER_46_501 VPWR VGND sg13g2_fill_2
XFILLER_15_965 VPWR VGND sg13g2_decap_8
XFILLER_30_913 VPWR VGND sg13g2_decap_8
XFILLER_42_784 VPWR VGND sg13g2_decap_8
XFILLER_41_261 VPWR VGND sg13g2_decap_4
XFILLER_6_663 VPWR VGND sg13g2_fill_2
XFILLER_6_652 VPWR VGND sg13g2_fill_1
XFILLER_5_151 VPWR VGND sg13g2_decap_8
X_4110_ _1046_ mydesign.pe_weights\[61\] mydesign.accum\[89\] _1071_ VPWR VGND sg13g2_a21o_1
X_5090_ _1931_ _1924_ _1933_ VPWR VGND sg13g2_xor2_1
XFILLER_25_1008 VPWR VGND sg13g2_decap_8
X_4041_ _0991_ VPWR _1014_ VGND _0990_ _0993_ sg13g2_o21ai_1
XFILLER_49_383 VPWR VGND sg13g2_decap_8
X_5992_ net142 VGND VPWR net953 mydesign.pe_weights\[30\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_4943_ mydesign.pe_weights\[38\] net528 mydesign.accum\[42\] _1799_ VPWR VGND sg13g2_nand3_1
XFILLER_21_902 VPWR VGND sg13g2_fill_1
X_4874_ _1749_ _1748_ _1750_ VPWR VGND sg13g2_xor2_1
XFILLER_21_946 VPWR VGND sg13g2_decap_8
X_3825_ VGND VPWR net572 _0816_ _0125_ _0817_ sg13g2_a21oi_1
X_3756_ _0763_ _0755_ _0760_ VPWR VGND sg13g2_nand2_1
X_5426_ _2236_ _2237_ _0306_ VPWR VGND sg13g2_nor2_1
X_3687_ _0690_ _0696_ _0697_ _0698_ VPWR VGND sg13g2_or3_1
XFILLER_0_817 VPWR VGND sg13g2_decap_8
X_5357_ mydesign.pe_inputs\[12\] net527 mydesign.accum\[19\] _2172_ VPWR VGND sg13g2_nand3_1
X_4308_ VGND VPWR net579 _1248_ _0176_ _1249_ sg13g2_a21oi_1
X_5288_ _2116_ _2113_ _2114_ VPWR VGND sg13g2_xnor2_1
X_4239_ _1184_ mydesign.accum\[81\] mydesign.pe_weights\[57\] net536 VPWR VGND sg13g2_and3_2
XFILLER_43_515 VPWR VGND sg13g2_decap_4
XFILLER_11_423 VPWR VGND sg13g2_fill_2
XFILLER_12_935 VPWR VGND sg13g2_decap_8
XFILLER_24_784 VPWR VGND sg13g2_fill_1
XFILLER_7_427 VPWR VGND sg13g2_decap_4
XFILLER_23_75 VPWR VGND sg13g2_fill_2
XFILLER_2_198 VPWR VGND sg13g2_fill_1
XFILLER_38_309 VPWR VGND sg13g2_fill_2
XFILLER_47_810 VPWR VGND sg13g2_decap_8
Xfanout491 net494 net491 VPWR VGND sg13g2_buf_8
Xfanout480 net482 net480 VPWR VGND sg13g2_buf_8
XFILLER_47_887 VPWR VGND sg13g2_decap_8
XFILLER_46_375 VPWR VGND sg13g2_fill_2
XFILLER_15_740 VPWR VGND sg13g2_fill_2
XFILLER_9_44 VPWR VGND sg13g2_fill_2
X_3610_ _0633_ _0629_ _0632_ VPWR VGND sg13g2_xnor2_1
X_4590_ mydesign.pe_inputs\[39\] mydesign.pe_weights\[51\] mydesign.accum\[70\] _1498_
+ VPWR VGND sg13g2_a21o_1
X_3541_ _0568_ _0545_ _0567_ VPWR VGND sg13g2_nand2_1
X_3472_ net627 VPWR _0508_ VGND net1086 net436 sg13g2_o21ai_1
X_5211_ _2043_ _2025_ _2041_ VPWR VGND sg13g2_xnor2_1
X_5142_ mydesign.pe_inputs\[23\] mydesign.pe_weights\[35\] mydesign.accum\[38\] _1982_
+ VPWR VGND sg13g2_a21o_1
XFILLER_38_821 VPWR VGND sg13g2_fill_1
X_5073_ _1917_ _1899_ _1916_ VPWR VGND sg13g2_nand2_1
X_4024_ _0998_ _0997_ _0987_ VPWR VGND sg13g2_nand2b_1
XFILLER_40_507 VPWR VGND sg13g2_decap_8
X_5975_ net207 VGND VPWR _0201_ mydesign.pe_weights\[33\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_4926_ VGND VPWR _2533_ net449 _0259_ _1784_ sg13g2_a21oi_1
XFILLER_33_581 VPWR VGND sg13g2_decap_4
X_4857_ _1732_ _1733_ _1734_ VPWR VGND sg13g2_nor2b_1
X_3808_ _0393_ _0801_ _0802_ _0803_ VPWR VGND sg13g2_nor3_2
X_4788_ _1668_ mydesign.pe_weights\[40\] mydesign.pe_inputs\[30\] VPWR VGND sg13g2_nand2_1
X_3739_ VGND VPWR mydesign.pe_inputs\[63\] _0658_ _0747_ mydesign.accum\[118\] sg13g2_a21oi_1
X_5409_ _2222_ _2202_ _2205_ _2221_ VPWR VGND sg13g2_and3_1
XFILLER_0_636 VPWR VGND sg13g2_decap_8
X_5849__71 VPWR VGND net71 sg13g2_tiehi
XFILLER_48_629 VPWR VGND sg13g2_decap_8
XFILLER_29_810 VPWR VGND sg13g2_fill_1
XFILLER_44_813 VPWR VGND sg13g2_decap_8
XFILLER_43_301 VPWR VGND sg13g2_decap_8
XFILLER_18_64 VPWR VGND sg13g2_fill_1
XFILLER_18_86 VPWR VGND sg13g2_decap_4
XFILLER_31_518 VPWR VGND sg13g2_fill_2
XFILLER_34_63 VPWR VGND sg13g2_decap_8
XFILLER_15_1007 VPWR VGND sg13g2_decap_8
Xheichips25_template_401 VPWR VGND uio_oe[2] sg13g2_tiehi
XFILLER_12_798 VPWR VGND sg13g2_fill_1
XFILLER_8_769 VPWR VGND sg13g2_fill_2
XFILLER_11_286 VPWR VGND sg13g2_decap_4
XFILLER_7_268 VPWR VGND sg13g2_fill_1
XFILLER_4_997 VPWR VGND sg13g2_decap_8
X_5855__63 VPWR VGND net63 sg13g2_tiehi
X_5870__33 VPWR VGND net33 sg13g2_tiehi
XFILLER_47_684 VPWR VGND sg13g2_decap_8
XFILLER_19_375 VPWR VGND sg13g2_fill_2
XFILLER_35_813 VPWR VGND sg13g2_fill_2
XFILLER_46_194 VPWR VGND sg13g2_decap_4
XFILLER_15_581 VPWR VGND sg13g2_decap_4
X_5760_ net615 VPWR _2510_ VGND _2591_ _1400_ sg13g2_o21ai_1
X_5691_ VGND VPWR net512 net457 _2471_ _2468_ sg13g2_a21oi_1
X_4711_ _1603_ _1595_ _1605_ VPWR VGND sg13g2_xor2_1
X_4642_ VGND VPWR _2550_ net437 _0218_ _1541_ sg13g2_a21oi_1
X_4573_ _1482_ _1480_ _1481_ VPWR VGND sg13g2_nand2_1
X_3524_ _0552_ _0534_ _0550_ VPWR VGND sg13g2_xnor2_1
X_3455_ _0495_ VPWR _0077_ VGND net602 _0492_ sg13g2_o21ai_1
X_3386_ VGND VPWR _0433_ _0434_ net514 mydesign.accum\[2\] sg13g2_a21oi_2
X_5125_ mydesign.pe_inputs\[23\] net530 mydesign.accum\[37\] _1966_ VPWR VGND sg13g2_a21o_1
X_5056_ _1899_ _1900_ _1901_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_673 VPWR VGND sg13g2_fill_2
X_4007_ _0964_ _0980_ _0981_ _0982_ VPWR VGND sg13g2_nor3_1
XFILLER_26_802 VPWR VGND sg13g2_decap_8
XFILLER_26_824 VPWR VGND sg13g2_fill_1
XFILLER_38_1007 VPWR VGND sg13g2_decap_8
X_5958_ net241 VGND VPWR _0184_ mydesign.pe_weights\[36\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_4909_ net612 VPWR _1776_ VGND net820 _1767_ sg13g2_o21ai_1
X_5889_ net374 VGND VPWR net708 mydesign.weights\[3\]\[7\] clknet_leaf_49_clk sg13g2_dfrbpq_1
XFILLER_1_901 VPWR VGND sg13g2_decap_8
XFILLER_0_400 VPWR VGND sg13g2_decap_8
XFILLER_49_916 VPWR VGND sg13g2_decap_8
XFILLER_1_978 VPWR VGND sg13g2_decap_8
XFILLER_0_488 VPWR VGND sg13g2_fill_1
Xhold41 mydesign.weights\[2\]\[9\] VPWR VGND net660 sg13g2_dlygate4sd3_1
Xhold30 mydesign.weights\[1\]\[19\] VPWR VGND net649 sg13g2_dlygate4sd3_1
XFILLER_48_437 VPWR VGND sg13g2_fill_1
Xhold52 mydesign.inputs\[3\]\[6\] VPWR VGND net671 sg13g2_dlygate4sd3_1
Xhold63 mydesign.inputs\[2\]\[17\] VPWR VGND net682 sg13g2_dlygate4sd3_1
Xhold74 mydesign.weights\[1\]\[21\] VPWR VGND net693 sg13g2_dlygate4sd3_1
XFILLER_29_85 VPWR VGND sg13g2_fill_2
Xhold85 mydesign.inputs\[2\]\[6\] VPWR VGND net704 sg13g2_dlygate4sd3_1
Xhold96 _0355_ VPWR VGND net715 sg13g2_dlygate4sd3_1
XFILLER_17_846 VPWR VGND sg13g2_decap_4
XFILLER_17_857 VPWR VGND sg13g2_fill_1
XFILLER_28_161 VPWR VGND sg13g2_fill_2
XFILLER_45_62 VPWR VGND sg13g2_decap_8
XFILLER_44_687 VPWR VGND sg13g2_decap_8
XFILLER_31_348 VPWR VGND sg13g2_fill_2
XFILLER_40_882 VPWR VGND sg13g2_decap_8
X_3240_ net608 net611 _2660_ VPWR VGND sg13g2_nor2_1
X_3171_ _2609_ VPWR _0001_ VGND net432 _2610_ sg13g2_o21ai_1
XFILLER_48_993 VPWR VGND sg13g2_decap_8
X_5812_ net130 VGND VPWR _0038_ mydesign.inputs\[1\]\[17\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5743_ _2501_ net748 _2500_ VPWR VGND sg13g2_nand2_1
X_6005__74 VPWR VGND net74 sg13g2_tiehi
XFILLER_31_860 VPWR VGND sg13g2_fill_1
X_5923__311 VPWR VGND net311 sg13g2_tiehi
X_5674_ VGND VPWR net409 _2459_ _0331_ _2460_ sg13g2_a21oi_1
X_4625_ mydesign.inputs\[2\]\[10\] mydesign.inputs\[2\]\[6\] net550 _1529_ VPWR VGND
+ sg13g2_mux2_1
X_4556_ _1466_ _1460_ _1465_ VPWR VGND sg13g2_nand2_1
XFILLER_2_709 VPWR VGND sg13g2_decap_4
X_3507_ net455 _0517_ net721 _0536_ VPWR VGND sg13g2_nand3_1
X_4487_ _1406_ net666 _1402_ VPWR VGND sg13g2_nand2_1
X_3438_ VGND VPWR _0412_ _0480_ _0481_ _2698_ sg13g2_a21oi_1
X_3369_ net513 mydesign.accum\[97\] mydesign.accum\[65\] mydesign.accum\[33\] mydesign.accum\[1\]
+ net506 _0418_ VPWR VGND sg13g2_mux4_1
XFILLER_46_908 VPWR VGND sg13g2_decap_8
X_5108_ _1950_ _1943_ _1949_ VPWR VGND sg13g2_nand2_1
Xheichips25_template_21 VPWR VGND uio_out[6] sg13g2_tielo
X_6088_ net380 VGND VPWR net1039 mydesign.accum\[10\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_5039_ VGND VPWR net583 _1888_ _0267_ _1889_ sg13g2_a21oi_1
XFILLER_15_54 VPWR VGND sg13g2_fill_2
XFILLER_22_871 VPWR VGND sg13g2_decap_8
XFILLER_5_547 VPWR VGND sg13g2_fill_1
XFILLER_5_536 VPWR VGND sg13g2_decap_4
Xoutput7 net7 uio_out[0] VPWR VGND sg13g2_buf_1
XFILLER_49_713 VPWR VGND sg13g2_decap_8
XFILLER_0_241 VPWR VGND sg13g2_decap_8
X_6078__88 VPWR VGND net88 sg13g2_tiehi
XFILLER_36_418 VPWR VGND sg13g2_fill_2
XFILLER_44_440 VPWR VGND sg13g2_fill_2
XFILLER_17_665 VPWR VGND sg13g2_decap_8
XFILLER_45_996 VPWR VGND sg13g2_decap_8
XFILLER_31_145 VPWR VGND sg13g2_fill_1
XFILLER_8_330 VPWR VGND sg13g2_decap_4
XFILLER_9_875 VPWR VGND sg13g2_decap_4
X_4410_ _1337_ _1313_ _1335_ VPWR VGND sg13g2_xnor2_1
X_5390_ _2183_ _2185_ _2203_ _2204_ VPWR VGND sg13g2_or3_1
X_4341_ net472 VPWR _1281_ VGND net579 net895 sg13g2_o21ai_1
X_4272_ mydesign.pe_inputs\[44\] net539 mydesign.accum\[83\] _1215_ VPWR VGND sg13g2_a21o_1
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
X_3223_ net1044 net842 _2647_ VPWR VGND sg13g2_and2_1
X_6011_ net46 VGND VPWR net893 mydesign.accum\[49\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_3154_ net555 net545 _2595_ VPWR VGND sg13g2_nor2b_2
XFILLER_48_790 VPWR VGND sg13g2_decap_8
X_6084__36 VPWR VGND net36 sg13g2_tiehi
XFILLER_27_418 VPWR VGND sg13g2_fill_2
X_3085_ VPWR _2526_ net939 VGND sg13g2_inv_1
XFILLER_36_930 VPWR VGND sg13g2_decap_8
XFILLER_35_462 VPWR VGND sg13g2_fill_1
XFILLER_35_473 VPWR VGND sg13g2_decap_8
X_3987_ VGND VPWR net564 _0961_ _0142_ _0962_ sg13g2_a21oi_1
XFILLER_10_307 VPWR VGND sg13g2_fill_2
X_5726_ _2491_ VPWR _0352_ VGND net604 _2490_ sg13g2_o21ai_1
X_5657_ _2431_ VPWR _2445_ VGND _2432_ _2433_ sg13g2_o21ai_1
XFILLER_11_1010 VPWR VGND sg13g2_decap_8
X_5588_ _2380_ _2375_ _2379_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_506 VPWR VGND sg13g2_fill_2
X_4608_ VGND VPWR net574 _1513_ _0211_ _1514_ sg13g2_a21oi_1
Xhold341 mydesign.accum\[117\] VPWR VGND net960 sg13g2_dlygate4sd3_1
X_4539_ _1448_ _1441_ _1450_ VPWR VGND sg13g2_xor2_1
Xhold352 mydesign.pe_weights\[53\] VPWR VGND net971 sg13g2_dlygate4sd3_1
Xhold330 mydesign.accum\[41\] VPWR VGND net949 sg13g2_dlygate4sd3_1
Xhold385 mydesign.accum\[127\] VPWR VGND net1004 sg13g2_dlygate4sd3_1
Xhold363 _0182_ VPWR VGND net982 sg13g2_dlygate4sd3_1
Xhold396 mydesign.pe_inputs\[57\] VPWR VGND net1015 sg13g2_dlygate4sd3_1
Xhold374 mydesign.pe_inputs\[43\] VPWR VGND net993 sg13g2_dlygate4sd3_1
XFILLER_46_705 VPWR VGND sg13g2_decap_8
XFILLER_27_941 VPWR VGND sg13g2_decap_8
XFILLER_14_613 VPWR VGND sg13g2_decap_4
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_42_933 VPWR VGND sg13g2_decap_8
XFILLER_26_484 VPWR VGND sg13g2_fill_2
XFILLER_9_105 VPWR VGND sg13g2_decap_4
XFILLER_10_830 VPWR VGND sg13g2_fill_1
XFILLER_5_311 VPWR VGND sg13g2_fill_1
XFILLER_6_867 VPWR VGND sg13g2_decap_8
XFILLER_47_9 VPWR VGND sg13g2_fill_1
XFILLER_49_521 VPWR VGND sg13g2_decap_8
XFILLER_49_510 VPWR VGND sg13g2_fill_1
XFILLER_49_554 VPWR VGND sg13g2_decap_8
XFILLER_49_587 VPWR VGND sg13g2_decap_8
XFILLER_18_974 VPWR VGND sg13g2_decap_8
XFILLER_45_793 VPWR VGND sg13g2_decap_8
X_4890_ _1763_ VPWR _0244_ VGND net603 _1761_ sg13g2_o21ai_1
X_3910_ _0883_ _0897_ _0898_ VPWR VGND sg13g2_nor2_1
X_3841_ net465 VPWR _0833_ VGND net572 net1010 sg13g2_o21ai_1
XFILLER_32_443 VPWR VGND sg13g2_decap_8
XFILLER_33_966 VPWR VGND sg13g2_decap_8
X_3772_ _0774_ VPWR _0115_ VGND net597 _0769_ sg13g2_o21ai_1
X_5511_ _2311_ VPWR _2313_ VGND _2291_ _2293_ sg13g2_o21ai_1
X_5442_ _2248_ net588 net521 mydesign.pe_weights\[20\] VPWR VGND sg13g2_and3_1
X_5373_ VGND VPWR net590 _2186_ _0303_ _2187_ sg13g2_a21oi_1
X_4324_ net579 VPWR _1265_ VGND _1263_ _1264_ sg13g2_o21ai_1
X_6020__386 VPWR VGND net386 sg13g2_tiehi
X_4255_ _1195_ _1198_ _1199_ VPWR VGND sg13g2_nor2_1
X_4186_ _1143_ mydesign.accum\[93\] _1142_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_1014 VPWR VGND sg13g2_decap_8
X_3206_ net616 _2633_ net692 _2636_ VPWR VGND sg13g2_nand3_1
X_3137_ VPWR _2578_ net808 VGND sg13g2_inv_1
XFILLER_42_229 VPWR VGND sg13g2_decap_8
X_6080__72 VPWR VGND net72 sg13g2_tiehi
X_5888__375 VPWR VGND net375 sg13g2_tiehi
XFILLER_24_988 VPWR VGND sg13g2_decap_8
XFILLER_10_137 VPWR VGND sg13g2_fill_1
X_5709_ mydesign.load_counter\[1\] _2605_ _2607_ _2483_ VPWR VGND sg13g2_nor3_1
XFILLER_3_837 VPWR VGND sg13g2_decap_4
Xhold160 mydesign.inputs\[1\]\[21\] VPWR VGND net779 sg13g2_dlygate4sd3_1
Xhold171 _0235_ VPWR VGND net790 sg13g2_dlygate4sd3_1
Xhold182 mydesign.inputs\[0\]\[19\] VPWR VGND net801 sg13g2_dlygate4sd3_1
Xhold193 _0217_ VPWR VGND net812 sg13g2_dlygate4sd3_1
X_5778__177 VPWR VGND net177 sg13g2_tiehi
Xfanout640 rst_n net640 VPWR VGND sg13g2_buf_8
XFILLER_46_568 VPWR VGND sg13g2_decap_4
XFILLER_18_259 VPWR VGND sg13g2_fill_1
XFILLER_27_771 VPWR VGND sg13g2_fill_1
XFILLER_15_944 VPWR VGND sg13g2_decap_8
XFILLER_42_774 VPWR VGND sg13g2_fill_1
XFILLER_42_752 VPWR VGND sg13g2_decap_8
X_6143__208 VPWR VGND net208 sg13g2_tiehi
XFILLER_18_1016 VPWR VGND sg13g2_decap_8
XFILLER_18_1027 VPWR VGND sg13g2_fill_2
XFILLER_26_292 VPWR VGND sg13g2_decap_4
XFILLER_41_284 VPWR VGND sg13g2_fill_1
XFILLER_30_969 VPWR VGND sg13g2_decap_8
XFILLER_2_870 VPWR VGND sg13g2_fill_1
XFILLER_49_340 VPWR VGND sg13g2_decap_8
X_4040_ _1012_ _1009_ _1013_ VPWR VGND sg13g2_xor2_1
X_5991_ net146 VGND VPWR net812 mydesign.pe_weights\[29\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_4942_ _1798_ mydesign.pe_weights\[37\] mydesign.pe_inputs\[25\] VPWR VGND sg13g2_nand2_1
X_4873_ VGND VPWR _1725_ _1733_ _1749_ _1732_ sg13g2_a21oi_1
XFILLER_21_925 VPWR VGND sg13g2_decap_8
X_3824_ net465 VPWR _0817_ VGND net572 net916 sg13g2_o21ai_1
X_3755_ _0761_ _0762_ _0110_ VPWR VGND sg13g2_nor2_1
X_3686_ VGND VPWR _0694_ _0695_ _0697_ _0674_ sg13g2_a21oi_1
X_5425_ net482 VPWR _2237_ VGND net590 net915 sg13g2_o21ai_1
X_5356_ _2171_ mydesign.pe_inputs\[13\] mydesign.pe_weights\[26\] VPWR VGND sg13g2_nand2_1
X_4307_ net471 VPWR _1249_ VGND net579 net933 sg13g2_o21ai_1
X_5287_ VPWR _2115_ _2114_ VGND sg13g2_inv_1
X_4238_ VGND VPWR net739 _1182_ _0172_ _1183_ sg13g2_a21oi_1
X_4169_ _1125_ _1123_ _1127_ VPWR VGND sg13g2_xor2_1
X_5931__295 VPWR VGND net295 sg13g2_tiehi
XFILLER_23_273 VPWR VGND sg13g2_fill_1
XFILLER_23_87 VPWR VGND sg13g2_fill_2
XFILLER_3_678 VPWR VGND sg13g2_fill_1
Xfanout492 net494 net492 VPWR VGND sg13g2_buf_8
Xfanout470 net472 net470 VPWR VGND sg13g2_buf_8
Xfanout481 net482 net481 VPWR VGND sg13g2_buf_8
XFILLER_47_866 VPWR VGND sg13g2_decap_8
XFILLER_34_505 VPWR VGND sg13g2_fill_1
XFILLER_42_593 VPWR VGND sg13g2_fill_1
XFILLER_9_56 VPWR VGND sg13g2_fill_2
X_5982__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_31_1013 VPWR VGND sg13g2_decap_8
X_3540_ _0567_ _0558_ _0565_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_995 VPWR VGND sg13g2_decap_8
X_3471_ VGND VPWR _2586_ _0506_ _0507_ net484 sg13g2_a21oi_1
X_5210_ _2042_ _2041_ _2025_ VPWR VGND sg13g2_nand2b_1
X_5141_ mydesign.pe_weights\[35\] mydesign.pe_inputs\[23\] mydesign.accum\[38\] _1981_
+ VPWR VGND sg13g2_nand3_1
X_5072_ _1916_ _1906_ _1915_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_811 VPWR VGND sg13g2_fill_2
XFILLER_38_800 VPWR VGND sg13g2_decap_8
X_4023_ _0996_ _0988_ _0997_ VPWR VGND sg13g2_xor2_1
XFILLER_49_170 VPWR VGND sg13g2_decap_8
XFILLER_38_855 VPWR VGND sg13g2_decap_4
XFILLER_37_310 VPWR VGND sg13g2_fill_1
XFILLER_38_888 VPWR VGND sg13g2_decap_8
X_5974_ net209 VGND VPWR net1034 mydesign.pe_weights\[32\] clknet_leaf_38_clk sg13g2_dfrbpq_2
XFILLER_40_519 VPWR VGND sg13g2_decap_8
X_4925_ net638 VPWR _1784_ VGND net1025 net449 sg13g2_o21ai_1
X_4856_ _1710_ _1731_ _1707_ _1733_ VPWR VGND sg13g2_nand3_1
XFILLER_20_221 VPWR VGND sg13g2_decap_4
XFILLER_21_744 VPWR VGND sg13g2_fill_1
X_3807_ mydesign.weights\[2\]\[15\] net550 _0802_ VPWR VGND sg13g2_nor2b_1
XFILLER_21_799 VPWR VGND sg13g2_fill_1
X_4787_ VGND VPWR net583 _1666_ _0237_ _1667_ sg13g2_a21oi_1
X_3738_ VGND VPWR net577 _0745_ _0109_ _0746_ sg13g2_a21oi_1
X_3669_ _0673_ _0680_ _0681_ VPWR VGND sg13g2_nor2b_1
XFILLER_47_1020 VPWR VGND sg13g2_decap_8
X_5408_ _2219_ _2198_ _2221_ VPWR VGND sg13g2_xor2_1
X_5339_ mydesign.pe_weights\[26\] net522 mydesign.accum\[18\] _2155_ VPWR VGND sg13g2_a21o_1
XFILLER_48_608 VPWR VGND sg13g2_decap_8
XFILLER_47_107 VPWR VGND sg13g2_fill_2
XFILLER_29_899 VPWR VGND sg13g2_decap_4
XFILLER_16_527 VPWR VGND sg13g2_fill_2
XFILLER_44_869 VPWR VGND sg13g2_decap_8
XFILLER_34_42 VPWR VGND sg13g2_decap_8
X_6066__194 VPWR VGND net194 sg13g2_tiehi
Xheichips25_template_402 VPWR VGND uio_oe[3] sg13g2_tiehi
XFILLER_34_75 VPWR VGND sg13g2_fill_2
XFILLER_7_203 VPWR VGND sg13g2_fill_2
XFILLER_4_976 VPWR VGND sg13g2_decap_8
X_6114__140 VPWR VGND net140 sg13g2_tiehi
XFILLER_22_8 VPWR VGND sg13g2_decap_8
XFILLER_38_129 VPWR VGND sg13g2_fill_2
XFILLER_47_663 VPWR VGND sg13g2_decap_8
XFILLER_34_313 VPWR VGND sg13g2_fill_1
XFILLER_22_519 VPWR VGND sg13g2_fill_2
X_5690_ _2466_ net834 _2470_ _0337_ VPWR VGND sg13g2_a21o_1
X_4710_ _1595_ _1603_ _1604_ VPWR VGND sg13g2_nor2_1
X_6045__278 VPWR VGND net278 sg13g2_tiehi
X_4641_ net625 VPWR _1541_ VGND mydesign.pe_weights\[30\] net437 sg13g2_o21ai_1
X_4572_ mydesign.pe_inputs\[38\] net537 mydesign.accum\[69\] _1481_ VPWR VGND sg13g2_a21o_1
XFILLER_6_280 VPWR VGND sg13g2_fill_1
X_3523_ _0551_ _0534_ _0550_ VPWR VGND sg13g2_nand2_1
X_3454_ _0495_ net425 _0493_ VPWR VGND sg13g2_nand2_1
XFILLER_41_0 VPWR VGND sg13g2_decap_8
X_3385_ net517 mydesign.accum\[34\] _0433_ VPWR VGND sg13g2_nor2b_1
X_5124_ net530 mydesign.pe_inputs\[23\] mydesign.accum\[37\] _1965_ VPWR VGND sg13g2_nand3_1
X_5055_ _1898_ VPWR _1900_ VGND _1896_ _1897_ sg13g2_o21ai_1
Xclkbuf_leaf_49_clk clknet_3_0__leaf_clk clknet_leaf_49_clk VPWR VGND sg13g2_buf_8
X_5891__371 VPWR VGND net371 sg13g2_tiehi
X_4006_ VGND VPWR _0978_ _0979_ _0981_ _0966_ sg13g2_a21oi_1
XFILLER_37_184 VPWR VGND sg13g2_fill_1
XFILLER_25_346 VPWR VGND sg13g2_fill_2
X_5957_ net243 VGND VPWR net994 mydesign.pe_inputs\[39\] clknet_leaf_40_clk sg13g2_dfrbpq_2
XFILLER_13_519 VPWR VGND sg13g2_fill_1
XFILLER_25_368 VPWR VGND sg13g2_fill_2
XFILLER_25_379 VPWR VGND sg13g2_fill_1
X_4908_ _1775_ net4 _1768_ VPWR VGND sg13g2_nand2_1
X_5888_ net375 VGND VPWR net702 mydesign.weights\[3\]\[6\] clknet_leaf_49_clk sg13g2_dfrbpq_1
XFILLER_21_585 VPWR VGND sg13g2_fill_1
X_4839_ _1715_ _1716_ _1717_ VPWR VGND sg13g2_and2_1
X_5781__173 VPWR VGND net173 sg13g2_tiehi
XFILLER_0_423 VPWR VGND sg13g2_decap_8
XFILLER_0_445 VPWR VGND sg13g2_decap_8
XFILLER_1_957 VPWR VGND sg13g2_decap_8
Xhold31 mydesign.inputs\[3\]\[10\] VPWR VGND net650 sg13g2_dlygate4sd3_1
Xhold20 _0077_ VPWR VGND net426 sg13g2_dlygate4sd3_1
Xhold53 mydesign.weights\[3\]\[5\] VPWR VGND net672 sg13g2_dlygate4sd3_1
Xhold42 _0293_ VPWR VGND net661 sg13g2_dlygate4sd3_1
Xhold64 mydesign.weights\[1\]\[16\] VPWR VGND net683 sg13g2_dlygate4sd3_1
Xhold86 mydesign.weights\[3\]\[2\] VPWR VGND net705 sg13g2_dlygate4sd3_1
Xhold75 mydesign.weights\[0\]\[22\] VPWR VGND net694 sg13g2_dlygate4sd3_1
Xhold97 mydesign.weights\[0\]\[25\] VPWR VGND net716 sg13g2_dlygate4sd3_1
XFILLER_21_1023 VPWR VGND sg13g2_decap_4
X_5852__67 VPWR VGND net67 sg13g2_tiehi
XFILLER_44_666 VPWR VGND sg13g2_decap_8
XFILLER_43_132 VPWR VGND sg13g2_decap_8
XFILLER_43_187 VPWR VGND sg13g2_decap_8
XFILLER_40_861 VPWR VGND sg13g2_decap_8
XFILLER_8_534 VPWR VGND sg13g2_fill_2
X_3170_ _2610_ net747 net618 VPWR VGND sg13g2_nand2_1
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_48_972 VPWR VGND sg13g2_decap_8
XFILLER_47_493 VPWR VGND sg13g2_fill_1
XFILLER_19_184 VPWR VGND sg13g2_fill_1
XFILLER_22_305 VPWR VGND sg13g2_fill_1
X_5811_ net131 VGND VPWR _0037_ mydesign.inputs\[1\]\[16\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5742_ net462 VPWR _2500_ VGND net608 _2663_ sg13g2_o21ai_1
X_5673_ net473 VPWR _2460_ VGND net409 _2459_ sg13g2_o21ai_1
XFILLER_31_894 VPWR VGND sg13g2_decap_8
X_4624_ VGND VPWR _2546_ net492 _0213_ _1528_ sg13g2_a21oi_1
X_4555_ _1464_ _1461_ _1465_ VPWR VGND sg13g2_xor2_1
X_3506_ _0533_ _0532_ _0535_ VPWR VGND sg13g2_xor2_1
X_4486_ _1405_ VPWR _0198_ VGND net599 _1401_ sg13g2_o21ai_1
X_3437_ net515 mydesign.accum\[111\] mydesign.accum\[79\] mydesign.accum\[47\] mydesign.accum\[15\]
+ net508 _0480_ VPWR VGND sg13g2_mux4_1
XFILLER_44_1023 VPWR VGND sg13g2_decap_4
X_3368_ VGND VPWR _0415_ _0416_ _0068_ _0417_ sg13g2_a21oi_1
X_5107_ _1947_ _1944_ _1949_ VPWR VGND sg13g2_xor2_1
X_3299_ _2632_ net605 net608 _2691_ VPWR VGND sg13g2_a21o_2
X_6087_ net388 VGND VPWR net929 mydesign.accum\[9\] clknet_leaf_34_clk sg13g2_dfrbpq_2
Xheichips25_template_22 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_26_611 VPWR VGND sg13g2_decap_4
X_5038_ net480 VPWR _1889_ VGND net583 net980 sg13g2_o21ai_1
XFILLER_41_636 VPWR VGND sg13g2_decap_8
XFILLER_21_371 VPWR VGND sg13g2_fill_2
XFILLER_21_382 VPWR VGND sg13g2_fill_1
XFILLER_31_76 VPWR VGND sg13g2_fill_1
Xoutput10 net10 uo_out[2] VPWR VGND sg13g2_buf_1
Xoutput8 net8 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_743 VPWR VGND sg13g2_fill_2
XFILLER_0_275 VPWR VGND sg13g2_fill_1
XFILLER_49_769 VPWR VGND sg13g2_decap_8
XFILLER_16_132 VPWR VGND sg13g2_decap_8
XFILLER_45_975 VPWR VGND sg13g2_decap_8
XFILLER_16_165 VPWR VGND sg13g2_decap_4
X_4340_ _1280_ _1279_ _1278_ VPWR VGND sg13g2_nand2b_1
X_4271_ net539 net536 mydesign.accum\[83\] _1214_ VPWR VGND sg13g2_nand3_1
X_3222_ _2646_ VPWR _0016_ VGND net598 _2641_ sg13g2_o21ai_1
X_6010_ net50 VGND VPWR net746 mydesign.accum\[48\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_3153_ VPWR _2594_ mydesign.inputs\[2\]\[7\] VGND sg13g2_inv_1
XFILLER_39_246 VPWR VGND sg13g2_fill_2
X_3084_ VPWR _2525_ net1000 VGND sg13g2_inv_1
XFILLER_36_986 VPWR VGND sg13g2_decap_8
XFILLER_23_625 VPWR VGND sg13g2_fill_1
X_3986_ net464 VPWR _0962_ VGND net565 net847 sg13g2_o21ai_1
X_5725_ net723 _2490_ net615 _2491_ VPWR VGND sg13g2_nand3_1
X_5656_ _2435_ VPWR _2444_ VGND _2429_ _2436_ sg13g2_o21ai_1
X_4607_ net473 VPWR _1514_ VGND net574 net843 sg13g2_o21ai_1
X_5587_ _2376_ _2378_ _2379_ VPWR VGND sg13g2_nor2_1
Xhold320 mydesign.pe_inputs\[14\] VPWR VGND net939 sg13g2_dlygate4sd3_1
Xhold342 mydesign.accum\[82\] VPWR VGND net961 sg13g2_dlygate4sd3_1
Xhold353 mydesign.accum\[116\] VPWR VGND net972 sg13g2_dlygate4sd3_1
X_4538_ _1441_ _1448_ _1449_ VPWR VGND sg13g2_nor2_1
Xhold331 _0261_ VPWR VGND net950 sg13g2_dlygate4sd3_1
Xhold364 mydesign.accum\[81\] VPWR VGND net983 sg13g2_dlygate4sd3_1
Xhold386 mydesign.accum\[37\] VPWR VGND net1005 sg13g2_dlygate4sd3_1
Xhold375 _0183_ VPWR VGND net994 sg13g2_dlygate4sd3_1
X_4469_ net480 VPWR _1393_ VGND net583 net909 sg13g2_o21ai_1
Xhold397 _0097_ VPWR VGND net1016 sg13g2_dlygate4sd3_1
X_6139_ net280 VGND VPWR net825 mydesign.weights\[3\]\[13\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_42_912 VPWR VGND sg13g2_decap_8
XFILLER_26_43 VPWR VGND sg13g2_fill_1
XFILLER_27_997 VPWR VGND sg13g2_decap_8
XFILLER_13_102 VPWR VGND sg13g2_fill_1
XFILLER_42_989 VPWR VGND sg13g2_decap_8
XFILLER_41_455 VPWR VGND sg13g2_fill_1
XFILLER_22_691 VPWR VGND sg13g2_decap_8
XFILLER_10_886 VPWR VGND sg13g2_decap_4
X_5941__275 VPWR VGND net275 sg13g2_tiehi
XFILLER_49_566 VPWR VGND sg13g2_fill_1
XFILLER_49_577 VPWR VGND sg13g2_fill_1
XFILLER_18_953 VPWR VGND sg13g2_decap_8
XFILLER_45_772 VPWR VGND sg13g2_decap_8
XFILLER_17_474 VPWR VGND sg13g2_fill_1
XFILLER_33_945 VPWR VGND sg13g2_decap_8
X_3840_ _0832_ _0815_ _0830_ VPWR VGND sg13g2_xnor2_1
X_3771_ _0774_ net707 _0770_ VPWR VGND sg13g2_nand2_1
XFILLER_9_651 VPWR VGND sg13g2_decap_8
X_5510_ _2291_ _2293_ _2311_ _2312_ VPWR VGND sg13g2_nor3_1
XFILLER_8_183 VPWR VGND sg13g2_decap_4
X_5441_ VGND VPWR _2521_ net445 _0311_ _2247_ sg13g2_a21oi_1
X_5372_ net481 VPWR _2187_ VGND net590 net992 sg13g2_o21ai_1
X_4323_ VGND VPWR _1244_ _1247_ _1264_ _1262_ sg13g2_a21oi_1
X_4254_ _1198_ _1196_ _1197_ VPWR VGND sg13g2_nand2_1
X_4185_ _1142_ mydesign.pe_weights\[63\] _1056_ VPWR VGND sg13g2_nand2_1
X_3205_ _2635_ VPWR _0010_ VGND _2519_ _2633_ sg13g2_o21ai_1
X_3136_ VPWR _2577_ net880 VGND sg13g2_inv_1
XFILLER_24_967 VPWR VGND sg13g2_decap_8
XFILLER_11_628 VPWR VGND sg13g2_fill_1
X_3969_ _0935_ mydesign.accum\[96\] _0944_ _0946_ VPWR VGND sg13g2_a21o_1
X_5708_ _2605_ _2639_ _2683_ _2482_ VPWR VGND sg13g2_nor3_1
X_5639_ _2419_ VPWR _2428_ VGND _2408_ _2420_ sg13g2_o21ai_1
XFILLER_3_816 VPWR VGND sg13g2_decap_8
Xhold150 mydesign.inputs\[1\]\[13\] VPWR VGND net769 sg13g2_dlygate4sd3_1
Xhold161 mydesign.inputs\[0\]\[16\] VPWR VGND net780 sg13g2_dlygate4sd3_1
Xhold172 mydesign.inputs\[1\]\[10\] VPWR VGND net791 sg13g2_dlygate4sd3_1
Xhold194 mydesign.pe_weights\[42\] VPWR VGND net813 sg13g2_dlygate4sd3_1
Xhold183 mydesign.weights\[1\]\[8\] VPWR VGND net802 sg13g2_dlygate4sd3_1
Xfanout630 net632 net630 VPWR VGND sg13g2_buf_8
XFILLER_46_525 VPWR VGND sg13g2_fill_2
XFILLER_2_1020 VPWR VGND sg13g2_decap_8
XFILLER_27_750 VPWR VGND sg13g2_decap_8
XFILLER_37_97 VPWR VGND sg13g2_fill_2
XFILLER_27_783 VPWR VGND sg13g2_decap_8
XFILLER_30_948 VPWR VGND sg13g2_decap_8
XFILLER_5_175 VPWR VGND sg13g2_decap_8
XFILLER_49_363 VPWR VGND sg13g2_fill_2
X_5990_ net166 VGND VPWR _0216_ mydesign.pe_weights\[28\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_4941_ _1797_ mydesign.pe_weights\[36\] mydesign.pe_inputs\[26\] VPWR VGND sg13g2_nand2_1
XFILLER_24_219 VPWR VGND sg13g2_fill_2
X_4872_ _1748_ _1747_ _1746_ VPWR VGND sg13g2_nand2b_1
X_3823_ _0814_ _0813_ _0816_ VPWR VGND sg13g2_xor2_1
X_3754_ net471 VPWR _0762_ VGND net570 net898 sg13g2_o21ai_1
XFILLER_9_481 VPWR VGND sg13g2_fill_1
X_3685_ _0696_ _0674_ _0694_ _0695_ VPWR VGND sg13g2_and3_1
X_5424_ VGND VPWR _2234_ _2235_ _2236_ net502 sg13g2_a21oi_1
X_5355_ _2170_ mydesign.pe_inputs\[14\] mydesign.pe_weights\[25\] VPWR VGND sg13g2_nand2_1
X_4306_ _1248_ _1247_ _1246_ VPWR VGND sg13g2_nand2b_1
X_5286_ _2097_ VPWR _2114_ VGND _2096_ _2099_ sg13g2_o21ai_1
X_4237_ net479 VPWR _1183_ VGND net739 _1182_ sg13g2_o21ai_1
X_4168_ _1123_ _1125_ _1126_ VPWR VGND sg13g2_nor2_1
XFILLER_28_536 VPWR VGND sg13g2_fill_2
XFILLER_43_506 VPWR VGND sg13g2_decap_4
X_3119_ VPWR _2560_ net993 VGND sg13g2_inv_1
X_4099_ net624 VPWR _1064_ VGND net811 net436 sg13g2_o21ai_1
XFILLER_43_528 VPWR VGND sg13g2_fill_1
Xfanout471 net472 net471 VPWR VGND sg13g2_buf_8
Xfanout482 net483 net482 VPWR VGND sg13g2_buf_8
Xfanout460 _0396_ net460 VPWR VGND sg13g2_buf_8
Xfanout493 net494 net493 VPWR VGND sg13g2_buf_8
XFILLER_47_845 VPWR VGND sg13g2_decap_8
XFILLER_46_377 VPWR VGND sg13g2_fill_1
XFILLER_14_241 VPWR VGND sg13g2_fill_2
XFILLER_9_46 VPWR VGND sg13g2_fill_1
XFILLER_7_974 VPWR VGND sg13g2_decap_8
X_3470_ _0505_ VPWR _0506_ VGND net544 _0504_ sg13g2_o21ai_1
X_5140_ _1980_ _1979_ _0277_ VPWR VGND sg13g2_nor2b_1
XFILLER_9_1026 VPWR VGND sg13g2_fill_2
X_5071_ _1912_ _1896_ _1915_ VPWR VGND sg13g2_xor2_1
X_4022_ _0996_ _0989_ _0994_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_834 VPWR VGND sg13g2_decap_8
X_5973_ net211 VGND VPWR _0199_ mydesign.inputs\[3\]\[15\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_4924_ VGND VPWR _2534_ net449 _0258_ _1783_ sg13g2_a21oi_1
X_5885__379 VPWR VGND net379 sg13g2_tiehi
X_4855_ VGND VPWR _1707_ _1710_ _1732_ _1731_ sg13g2_a21oi_1
X_3806_ net550 mydesign.weights\[2\]\[19\] _0801_ VPWR VGND sg13g2_nor2_1
XFILLER_21_767 VPWR VGND sg13g2_fill_2
X_4786_ net480 VPWR _1667_ VGND net583 net892 sg13g2_o21ai_1
X_3737_ net471 VPWR _0746_ VGND net580 net960 sg13g2_o21ai_1
X_3668_ _0680_ _0663_ _0679_ VPWR VGND sg13g2_xnor2_1
X_3599_ _0623_ _0622_ _0608_ VPWR VGND sg13g2_nand2b_1
X_5407_ _2198_ _2219_ _2220_ VPWR VGND sg13g2_nor2b_1
X_5338_ net522 mydesign.pe_weights\[26\] mydesign.accum\[18\] _2154_ VPWR VGND sg13g2_nand3_1
X_5269_ _2015_ mydesign.pe_weights\[31\] mydesign.accum\[29\] _2098_ VPWR VGND sg13g2_a21o_1
XFILLER_16_506 VPWR VGND sg13g2_decap_4
XFILLER_44_848 VPWR VGND sg13g2_decap_8
XFILLER_16_539 VPWR VGND sg13g2_fill_1
XFILLER_24_572 VPWR VGND sg13g2_decap_8
Xheichips25_template_403 VPWR VGND uio_oe[4] sg13g2_tiehi
XFILLER_4_955 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_fill_2
XFILLER_3_498 VPWR VGND sg13g2_fill_2
X_6073__144 VPWR VGND net144 sg13g2_tiehi
XFILLER_19_300 VPWR VGND sg13g2_fill_1
XFILLER_47_642 VPWR VGND sg13g2_decap_8
XFILLER_19_333 VPWR VGND sg13g2_fill_1
XFILLER_35_815 VPWR VGND sg13g2_fill_1
X_5830__109 VPWR VGND net109 sg13g2_tiehi
XFILLER_34_303 VPWR VGND sg13g2_fill_2
XFILLER_30_564 VPWR VGND sg13g2_decap_4
X_4640_ VGND VPWR _2551_ net437 _0217_ _1540_ sg13g2_a21oi_1
X_4571_ net537 mydesign.pe_inputs\[38\] mydesign.accum\[69\] _1480_ VPWR VGND sg13g2_nand3_1
X_3522_ _0550_ _0540_ _0548_ VPWR VGND sg13g2_xnor2_1
X_3453_ _0494_ VPWR _0076_ VGND net604 _0492_ sg13g2_o21ai_1
X_3384_ mydesign.accum\[98\] mydesign.accum\[66\] net512 _0432_ VPWR VGND sg13g2_mux2_1
X_5123_ _1964_ mydesign.pe_weights\[35\] mydesign.pe_inputs\[22\] VPWR VGND sg13g2_nand2_1
X_5054_ _1896_ _1897_ _1898_ _1899_ VPWR VGND sg13g2_nor3_1
XFILLER_38_642 VPWR VGND sg13g2_decap_4
X_4005_ _0980_ _0966_ _0978_ _0979_ VPWR VGND sg13g2_and3_1
XFILLER_38_675 VPWR VGND sg13g2_fill_1
X_5956_ net245 VGND VPWR net982 mydesign.pe_inputs\[38\] clknet_leaf_40_clk sg13g2_dfrbpq_2
X_4907_ VGND VPWR _1767_ _1773_ _0250_ net854 sg13g2_a21oi_1
X_5887_ net376 VGND VPWR net673 mydesign.weights\[3\]\[5\] clknet_leaf_49_clk sg13g2_dfrbpq_1
XFILLER_21_531 VPWR VGND sg13g2_fill_1
X_4838_ _1692_ _1694_ _1714_ _1716_ VPWR VGND sg13g2_or3_1
X_4769_ VGND VPWR _2543_ net451 _0233_ _1653_ sg13g2_a21oi_1
XFILLER_1_936 VPWR VGND sg13g2_decap_8
Xhold10 mydesign.inputs\[3\]\[8\] VPWR VGND net416 sg13g2_dlygate4sd3_1
Xhold32 _0322_ VPWR VGND net651 sg13g2_dlygate4sd3_1
XFILLER_0_479 VPWR VGND sg13g2_decap_8
Xhold21 mydesign.weights\[2\]\[10\] VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold54 _0113_ VPWR VGND net673 sg13g2_dlygate4sd3_1
Xhold65 mydesign.accum\[72\] VPWR VGND net684 sg13g2_dlygate4sd3_1
Xhold43 mydesign.weights\[2\]\[19\] VPWR VGND net662 sg13g2_dlygate4sd3_1
XFILLER_21_1002 VPWR VGND sg13g2_decap_8
Xhold98 mydesign.weights\[3\]\[1\] VPWR VGND net717 sg13g2_dlygate4sd3_1
Xhold87 _0342_ VPWR VGND net706 sg13g2_dlygate4sd3_1
Xhold76 mydesign.weights\[2\]\[8\] VPWR VGND net695 sg13g2_dlygate4sd3_1
XFILLER_45_31 VPWR VGND sg13g2_decap_4
XFILLER_28_163 VPWR VGND sg13g2_fill_1
XFILLER_29_675 VPWR VGND sg13g2_fill_2
XFILLER_44_645 VPWR VGND sg13g2_decap_8
XFILLER_16_369 VPWR VGND sg13g2_fill_2
XFILLER_8_568 VPWR VGND sg13g2_decap_4
XFILLER_6_1007 VPWR VGND sg13g2_decap_8
XFILLER_48_951 VPWR VGND sg13g2_decap_8
X_5951__255 VPWR VGND net255 sg13g2_tiehi
X_5810_ net133 VGND VPWR _0036_ mydesign.inputs\[2\]\[19\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_16_881 VPWR VGND sg13g2_fill_1
X_5741_ _2499_ VPWR _0359_ VGND net598 _2495_ sg13g2_o21ai_1
X_5672_ VGND VPWR _2458_ _2459_ _2457_ _2456_ sg13g2_a21oi_2
X_4623_ net625 VPWR _1528_ VGND net489 _1527_ sg13g2_o21ai_1
X_4554_ _1464_ _1462_ _1463_ VPWR VGND sg13g2_nand2_1
X_3505_ _0532_ _0533_ _0534_ VPWR VGND sg13g2_nor2_1
X_4485_ _1405_ net422 _1402_ VPWR VGND sg13g2_nand2_1
XFILLER_44_1002 VPWR VGND sg13g2_decap_8
X_3436_ VGND VPWR _0470_ _0478_ _0074_ _0479_ sg13g2_a21oi_1
X_3367_ net623 VPWR _0417_ VGND net1081 net430 sg13g2_o21ai_1
X_5106_ VGND VPWR _1948_ _1947_ _1944_ sg13g2_or2_1
X_6086_ net396 VGND VPWR net730 mydesign.accum\[8\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3298_ _2670_ net787 _2690_ _0048_ VPWR VGND sg13g2_mux2_1
X_5037_ _1888_ _1884_ _1887_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_984 VPWR VGND sg13g2_decap_8
XFILLER_15_56 VPWR VGND sg13g2_fill_1
X_5939_ net279 VGND VPWR _0165_ mydesign.pe_inputs\[41\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_22_895 VPWR VGND sg13g2_decap_4
X_6011__46 VPWR VGND net46 sg13g2_tiehi
Xoutput9 net9 uo_out[1] VPWR VGND sg13g2_buf_1
Xoutput11 net11 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_722 VPWR VGND sg13g2_fill_1
XFILLER_49_748 VPWR VGND sg13g2_decap_8
XFILLER_29_450 VPWR VGND sg13g2_decap_4
XFILLER_45_954 VPWR VGND sg13g2_decap_8
XFILLER_16_122 VPWR VGND sg13g2_decap_4
XFILLER_31_103 VPWR VGND sg13g2_decap_4
X_5829__111 VPWR VGND net111 sg13g2_tiehi
XFILLER_13_895 VPWR VGND sg13g2_fill_1
X_4270_ _1213_ mydesign.pe_weights\[58\] mydesign.pe_inputs\[45\] VPWR VGND sg13g2_nand2_1
X_5979__199 VPWR VGND net199 sg13g2_tiehi
XFILLER_28_1019 VPWR VGND sg13g2_decap_8
X_3221_ _2646_ net642 _2642_ VPWR VGND sg13g2_nand2_1
XFILLER_39_214 VPWR VGND sg13g2_fill_2
X_3152_ VPWR _2593_ net411 VGND sg13g2_inv_1
X_3083_ VPWR _2524_ net521 VGND sg13g2_inv_1
XFILLER_36_965 VPWR VGND sg13g2_decap_8
X_3985_ _0961_ _0945_ _0960_ VPWR VGND sg13g2_xnor2_1
X_5724_ _2619_ _2621_ net611 _2490_ VPWR VGND sg13g2_nand3_1
XFILLER_31_681 VPWR VGND sg13g2_decap_4
X_5655_ VGND VPWR net586 _2442_ _0329_ _2443_ sg13g2_a21oi_1
X_4606_ _1513_ _1509_ _1512_ VPWR VGND sg13g2_xnor2_1
X_6001__90 VPWR VGND net90 sg13g2_tiehi
X_5586_ VGND VPWR mydesign.pe_inputs\[6\] net523 _2378_ mydesign.accum\[2\] sg13g2_a21oi_1
Xhold310 _0313_ VPWR VGND net929 sg13g2_dlygate4sd3_1
Xhold332 mydesign.accum\[85\] VPWR VGND net951 sg13g2_dlygate4sd3_1
Xhold343 _0174_ VPWR VGND net962 sg13g2_dlygate4sd3_1
X_4537_ _1446_ _1425_ _1448_ VPWR VGND sg13g2_xor2_1
Xhold321 mydesign.accum\[103\] VPWR VGND net940 sg13g2_dlygate4sd3_1
Xhold376 mydesign.pe_weights\[56\] VPWR VGND net995 sg13g2_dlygate4sd3_1
Xhold365 _0173_ VPWR VGND net984 sg13g2_dlygate4sd3_1
Xhold354 mydesign.accum\[119\] VPWR VGND net973 sg13g2_dlygate4sd3_1
Xhold387 mydesign.accum\[100\] VPWR VGND net1006 sg13g2_dlygate4sd3_1
X_4468_ VGND VPWR _1390_ _1391_ _1392_ net502 sg13g2_a21oi_1
Xhold398 mydesign.pe_weights\[18\] VPWR VGND net1017 sg13g2_dlygate4sd3_1
X_3419_ net515 mydesign.accum\[109\] mydesign.accum\[77\] mydesign.accum\[45\] mydesign.accum\[13\]
+ net508 _0464_ VPWR VGND sg13g2_mux4_1
X_6138_ net296 VGND VPWR net987 mydesign.weights\[3\]\[12\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4399_ _1326_ mydesign.pe_weights\[53\] mydesign.pe_inputs\[42\] VPWR VGND sg13g2_nand2_1
X_6069_ net188 VGND VPWR net657 mydesign.weights\[2\]\[11\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_27_976 VPWR VGND sg13g2_decap_8
XFILLER_41_423 VPWR VGND sg13g2_decap_8
XFILLER_26_88 VPWR VGND sg13g2_decap_8
XFILLER_26_99 VPWR VGND sg13g2_fill_2
XFILLER_42_968 VPWR VGND sg13g2_decap_8
XFILLER_13_169 VPWR VGND sg13g2_fill_2
XFILLER_10_854 VPWR VGND sg13g2_decap_8
XFILLER_42_98 VPWR VGND sg13g2_decap_4
X_5906__341 VPWR VGND net341 sg13g2_tiehi
XFILLER_6_847 VPWR VGND sg13g2_fill_2
XFILLER_45_751 VPWR VGND sg13g2_decap_8
XFILLER_33_924 VPWR VGND sg13g2_decap_8
XFILLER_44_294 VPWR VGND sg13g2_fill_2
XFILLER_32_456 VPWR VGND sg13g2_fill_2
X_3770_ _0773_ VPWR _0114_ VGND net599 _0769_ sg13g2_o21ai_1
XFILLER_13_670 VPWR VGND sg13g2_fill_2
XFILLER_34_1012 VPWR VGND sg13g2_decap_8
X_5440_ net635 VPWR _2247_ VGND net946 net444 sg13g2_o21ai_1
X_5371_ _2184_ _2167_ _2186_ VPWR VGND sg13g2_xor2_1
X_4322_ _1263_ _1244_ _1247_ _1262_ VPWR VGND sg13g2_and3_1
X_5803__147 VPWR VGND net147 sg13g2_tiehi
X_4253_ net536 mydesign.pe_weights\[58\] mydesign.accum\[82\] _1197_ VPWR VGND sg13g2_a21o_1
X_3204_ net616 _2633_ net675 _2635_ VPWR VGND sg13g2_nand3_1
X_4184_ _1141_ mydesign.pe_weights\[62\] _1061_ VPWR VGND sg13g2_nand2_1
X_3135_ VPWR _2576_ net838 VGND sg13g2_inv_1
XFILLER_27_239 VPWR VGND sg13g2_fill_2
XFILLER_24_946 VPWR VGND sg13g2_decap_8
X_3968_ _0935_ _0944_ mydesign.accum\[96\] _0945_ VPWR VGND sg13g2_nand3_1
X_5707_ _2354_ net610 net609 _2481_ VPWR VGND sg13g2_a21o_2
X_3899_ VGND VPWR _0888_ _0887_ _0868_ sg13g2_or2_1
X_5638_ _2423_ VPWR _2427_ VGND _2404_ _2424_ sg13g2_o21ai_1
X_5569_ VGND VPWR net749 _2361_ _0324_ _2362_ sg13g2_a21oi_1
Xhold162 mydesign.weights\[0\]\[15\] VPWR VGND net781 sg13g2_dlygate4sd3_1
Xhold151 mydesign.weights\[1\]\[10\] VPWR VGND net770 sg13g2_dlygate4sd3_1
Xhold140 _0300_ VPWR VGND net759 sg13g2_dlygate4sd3_1
Xhold173 mydesign.inputs\[0\]\[23\] VPWR VGND net792 sg13g2_dlygate4sd3_1
Xhold184 mydesign.weights\[0\]\[13\] VPWR VGND net803 sg13g2_dlygate4sd3_1
Xhold195 _0234_ VPWR VGND net814 sg13g2_dlygate4sd3_1
Xfanout631 net632 net631 VPWR VGND sg13g2_buf_8
Xfanout620 net621 net620 VPWR VGND sg13g2_buf_8
XFILLER_26_250 VPWR VGND sg13g2_fill_2
XFILLER_15_979 VPWR VGND sg13g2_decap_8
XFILLER_42_798 VPWR VGND sg13g2_decap_8
XFILLER_30_927 VPWR VGND sg13g2_decap_8
XFILLER_10_662 VPWR VGND sg13g2_fill_2
XFILLER_10_684 VPWR VGND sg13g2_decap_4
XFILLER_5_165 VPWR VGND sg13g2_fill_1
XFILLER_49_320 VPWR VGND sg13g2_decap_8
XFILLER_1_382 VPWR VGND sg13g2_fill_1
XFILLER_37_504 VPWR VGND sg13g2_decap_8
XFILLER_49_397 VPWR VGND sg13g2_decap_8
X_4940_ VGND VPWR net585 _1795_ _0261_ _1796_ sg13g2_a21oi_1
X_4871_ _1730_ _1745_ _1727_ _1747_ VPWR VGND sg13g2_nand3_1
X_6048__266 VPWR VGND net266 sg13g2_tiehi
X_3822_ mydesign.pe_inputs\[56\] _0783_ net688 _0815_ VPWR VGND _0813_ sg13g2_nand4_1
XFILLER_32_264 VPWR VGND sg13g2_decap_4
X_6541_ mydesign.valid_out net7 VPWR VGND sg13g2_buf_1
X_3753_ VGND VPWR _0759_ _0760_ _0761_ net502 sg13g2_a21oi_1
X_3684_ _0691_ VPWR _0695_ VGND _0692_ _0693_ sg13g2_o21ai_1
X_5423_ _2233_ VPWR _2235_ VGND _2220_ _2223_ sg13g2_o21ai_1
X_5354_ _2169_ mydesign.pe_inputs\[15\] mydesign.pe_weights\[24\] VPWR VGND sg13g2_nand2_1
X_4305_ _1245_ VPWR _1247_ VGND _1225_ _1227_ sg13g2_o21ai_1
X_5285_ _2113_ _2112_ _2111_ VPWR VGND sg13g2_nand2b_1
X_4236_ net502 _2567_ _2571_ _1182_ VPWR VGND sg13g2_nor3_1
X_4167_ _1125_ mydesign.accum\[92\] _1124_ VPWR VGND sg13g2_xnor2_1
X_3118_ _2559_ net910 VPWR VGND sg13g2_inv_2
X_4098_ VGND VPWR _2578_ net436 _0152_ _1063_ sg13g2_a21oi_1
XFILLER_24_732 VPWR VGND sg13g2_decap_8
XFILLER_12_916 VPWR VGND sg13g2_fill_1
XFILLER_24_776 VPWR VGND sg13g2_fill_2
XFILLER_12_949 VPWR VGND sg13g2_decap_8
X_6142__232 VPWR VGND net232 sg13g2_tiehi
XFILLER_20_982 VPWR VGND sg13g2_decap_8
XFILLER_23_89 VPWR VGND sg13g2_fill_1
Xfanout450 net451 net450 VPWR VGND sg13g2_buf_8
XFILLER_47_824 VPWR VGND sg13g2_decap_8
Xfanout461 _0390_ net461 VPWR VGND sg13g2_buf_8
Xfanout483 _2660_ net483 VPWR VGND sg13g2_buf_8
Xfanout472 net483 net472 VPWR VGND sg13g2_buf_8
XFILLER_46_312 VPWR VGND sg13g2_fill_2
XFILLER_19_526 VPWR VGND sg13g2_fill_2
XFILLER_19_548 VPWR VGND sg13g2_decap_4
Xfanout494 _2602_ net494 VPWR VGND sg13g2_buf_8
X_5910__337 VPWR VGND net337 sg13g2_tiehi
XFILLER_15_787 VPWR VGND sg13g2_fill_2
XFILLER_14_275 VPWR VGND sg13g2_fill_1
XFILLER_14_286 VPWR VGND sg13g2_fill_2
XFILLER_10_470 VPWR VGND sg13g2_fill_2
XFILLER_11_982 VPWR VGND sg13g2_decap_8
XFILLER_9_1005 VPWR VGND sg13g2_decap_8
XFILLER_36_4 VPWR VGND sg13g2_fill_1
X_5070_ _1896_ _1912_ _1914_ VPWR VGND sg13g2_nor2_1
XFILLER_2_691 VPWR VGND sg13g2_fill_1
X_6019__390 VPWR VGND net390 sg13g2_tiehi
X_4021_ _0995_ _0989_ _0994_ VPWR VGND sg13g2_nand2_1
XFILLER_37_301 VPWR VGND sg13g2_decap_8
XFILLER_37_334 VPWR VGND sg13g2_fill_2
X_5972_ net213 VGND VPWR _0198_ mydesign.inputs\[3\]\[14\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_4923_ net638 VPWR _1783_ VGND net525 net449 sg13g2_o21ai_1
X_4854_ _1731_ _1726_ _1729_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_735 VPWR VGND sg13g2_decap_8
X_3805_ _0397_ _0798_ _0799_ _0800_ VPWR VGND sg13g2_nor3_1
X_4785_ _1664_ _1663_ _1666_ VPWR VGND sg13g2_xor2_1
X_3736_ _0745_ _0730_ _0744_ VPWR VGND sg13g2_xnor2_1
X_5961__235 VPWR VGND net235 sg13g2_tiehi
X_6102__260 VPWR VGND net260 sg13g2_tiehi
X_3667_ _0679_ _0676_ _0677_ VPWR VGND sg13g2_xnor2_1
X_3598_ _0620_ _0606_ _0622_ VPWR VGND sg13g2_xor2_1
X_5406_ _2217_ _2216_ _2219_ VPWR VGND sg13g2_xor2_1
XFILLER_0_606 VPWR VGND sg13g2_decap_8
X_5337_ _2153_ mydesign.pe_inputs\[13\] mydesign.pe_weights\[25\] VPWR VGND sg13g2_nand2_1
X_5268_ mydesign.pe_weights\[31\] _2015_ mydesign.accum\[29\] _2097_ VPWR VGND sg13g2_nand3_1
X_4219_ VGND VPWR net569 _1172_ _0163_ _1173_ sg13g2_a21oi_1
XFILLER_18_12 VPWR VGND sg13g2_fill_2
XFILLER_18_23 VPWR VGND sg13g2_fill_2
X_5199_ VGND VPWR mydesign.accum\[24\] _2022_ _2032_ _2030_ sg13g2_a21oi_1
XFILLER_29_824 VPWR VGND sg13g2_decap_8
XFILLER_28_334 VPWR VGND sg13g2_fill_2
XFILLER_29_868 VPWR VGND sg13g2_decap_8
XFILLER_44_827 VPWR VGND sg13g2_decap_8
XFILLER_43_315 VPWR VGND sg13g2_fill_1
XFILLER_43_359 VPWR VGND sg13g2_fill_2
Xheichips25_template_404 VPWR VGND uio_oe[5] sg13g2_tiehi
XFILLER_34_77 VPWR VGND sg13g2_fill_1
XFILLER_7_205 VPWR VGND sg13g2_fill_1
XFILLER_11_256 VPWR VGND sg13g2_fill_2
XFILLER_3_411 VPWR VGND sg13g2_fill_2
XFILLER_3_444 VPWR VGND sg13g2_fill_1
XFILLER_3_433 VPWR VGND sg13g2_decap_8
XFILLER_47_621 VPWR VGND sg13g2_decap_8
XFILLER_47_698 VPWR VGND sg13g2_decap_8
XFILLER_43_893 VPWR VGND sg13g2_decap_8
XFILLER_42_392 VPWR VGND sg13g2_fill_2
XFILLER_30_543 VPWR VGND sg13g2_decap_8
X_4570_ _1479_ mydesign.pe_weights\[50\] mydesign.pe_inputs\[39\] VPWR VGND sg13g2_nand2_1
X_3521_ _0549_ _0548_ _0540_ VPWR VGND sg13g2_nand2b_1
X_3452_ _0494_ net414 _0493_ VPWR VGND sg13g2_nand2_1
X_3383_ net515 mydesign.accum\[114\] mydesign.accum\[82\] mydesign.accum\[50\] mydesign.accum\[18\]
+ net509 _0431_ VPWR VGND sg13g2_mux4_1
X_5122_ _1950_ VPWR _1963_ VGND _1942_ _1951_ sg13g2_o21ai_1
X_5053_ _1898_ mydesign.pe_weights\[32\] mydesign.pe_inputs\[21\] VPWR VGND sg13g2_nand2_1
X_5846__77 VPWR VGND net77 sg13g2_tiehi
X_4004_ _0976_ _0975_ _0953_ _0979_ VPWR VGND sg13g2_a21o_1
XFILLER_41_808 VPWR VGND sg13g2_fill_2
X_5955_ net247 VGND VPWR _0181_ mydesign.pe_inputs\[37\] clknet_leaf_44_clk sg13g2_dfrbpq_2
X_4906_ net613 VPWR _1774_ VGND net853 _1767_ sg13g2_o21ai_1
X_5886_ net377 VGND VPWR net412 mydesign.weights\[3\]\[4\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_34_893 VPWR VGND sg13g2_decap_8
XFILLER_21_554 VPWR VGND sg13g2_fill_1
XFILLER_33_392 VPWR VGND sg13g2_fill_2
X_4837_ _1714_ VPWR _1715_ VGND _1692_ _1694_ sg13g2_o21ai_1
X_4768_ net637 VPWR _1653_ VGND mydesign.pe_weights\[25\] net451 sg13g2_o21ai_1
X_4699_ _1589_ VPWR _1593_ VGND _1571_ _1590_ sg13g2_o21ai_1
X_3719_ net470 VPWR _0729_ VGND net577 net972 sg13g2_o21ai_1
XFILLER_1_915 VPWR VGND sg13g2_decap_8
XFILLER_0_414 VPWR VGND sg13g2_fill_1
Xhold11 _0320_ VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold22 _0294_ VPWR VGND net641 sg13g2_dlygate4sd3_1
Xhold44 _0012_ VPWR VGND net663 sg13g2_dlygate4sd3_1
Xhold33 mydesign.inputs\[2\]\[15\] VPWR VGND net652 sg13g2_dlygate4sd3_1
XFILLER_29_77 VPWR VGND sg13g2_fill_2
XFILLER_29_621 VPWR VGND sg13g2_fill_1
Xhold55 mydesign.weights\[1\]\[23\] VPWR VGND net674 sg13g2_dlygate4sd3_1
Xhold88 mydesign.weights\[3\]\[7\] VPWR VGND net707 sg13g2_dlygate4sd3_1
Xhold99 _0341_ VPWR VGND net718 sg13g2_dlygate4sd3_1
Xhold66 _0188_ VPWR VGND net685 sg13g2_dlygate4sd3_1
Xhold77 _0292_ VPWR VGND net696 sg13g2_dlygate4sd3_1
XFILLER_16_304 VPWR VGND sg13g2_fill_2
XFILLER_17_816 VPWR VGND sg13g2_decap_4
XFILLER_16_348 VPWR VGND sg13g2_decap_4
XFILLER_43_167 VPWR VGND sg13g2_decap_8
XFILLER_32_819 VPWR VGND sg13g2_decap_8
XFILLER_40_896 VPWR VGND sg13g2_decap_8
XFILLER_4_753 VPWR VGND sg13g2_fill_1
XFILLER_4_786 VPWR VGND sg13g2_fill_2
XFILLER_4_775 VPWR VGND sg13g2_fill_2
XFILLER_4_764 VPWR VGND sg13g2_decap_8
XFILLER_48_930 VPWR VGND sg13g2_decap_8
XFILLER_0_992 VPWR VGND sg13g2_decap_8
XFILLER_19_142 VPWR VGND sg13g2_fill_1
XFILLER_35_657 VPWR VGND sg13g2_fill_2
X_5740_ _2499_ net722 _2495_ VPWR VGND sg13g2_nand2_1
X_5671_ net587 VPWR _2458_ VGND _2456_ _2457_ sg13g2_o21ai_1
X_4622_ _1524_ VPWR _1527_ VGND _1525_ _1526_ sg13g2_o21ai_1
X_4553_ mydesign.pe_inputs\[37\] net537 mydesign.accum\[68\] _1463_ VPWR VGND sg13g2_a21o_1
X_4484_ _1404_ VPWR _0197_ VGND net601 _1401_ sg13g2_o21ai_1
X_3504_ _0533_ _0501_ _0517_ VPWR VGND sg13g2_nand2_1
X_3435_ net622 VPWR _0479_ VGND net1072 net430 sg13g2_o21ai_1
X_3366_ VPWR VGND _0406_ _0414_ _0405_ net458 _0416_ _0404_ sg13g2_a221oi_1
X_3297_ _2669_ net772 _2690_ _0047_ VPWR VGND sg13g2_mux2_1
X_5105_ _1947_ _1945_ _1946_ VPWR VGND sg13g2_nand2_1
X_6085_ net28 VGND VPWR net947 mydesign.pe_inputs\[7\] clknet_leaf_35_clk sg13g2_dfrbpq_1
XFILLER_39_963 VPWR VGND sg13g2_decap_8
X_5036_ _1887_ _1885_ _1886_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_602 VPWR VGND sg13g2_fill_1
X_5938_ net281 VGND VPWR net1051 mydesign.pe_inputs\[40\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_22_863 VPWR VGND sg13g2_fill_2
X_5869_ net35 VGND VPWR _0095_ mydesign.accum\[127\] clknet_leaf_17_clk sg13g2_dfrbpq_2
Xoutput12 net12 uo_out[4] VPWR VGND sg13g2_buf_1
X_5898__357 VPWR VGND net357 sg13g2_tiehi
XFILLER_0_255 VPWR VGND sg13g2_decap_4
XFILLER_49_727 VPWR VGND sg13g2_decap_8
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_45_933 VPWR VGND sg13g2_decap_8
XFILLER_44_410 VPWR VGND sg13g2_decap_8
XFILLER_17_679 VPWR VGND sg13g2_decap_8
XFILLER_13_874 VPWR VGND sg13g2_fill_1
XFILLER_4_550 VPWR VGND sg13g2_decap_4
X_3220_ _2645_ VPWR _0015_ VGND net600 _2641_ sg13g2_o21ai_1
X_3151_ VPWR _2592_ mydesign.weights\[0\]\[24\] VGND sg13g2_inv_1
XFILLER_39_248 VPWR VGND sg13g2_fill_1
X_3082_ VPWR _2523_ net934 VGND sg13g2_inv_1
XFILLER_35_432 VPWR VGND sg13g2_fill_1
XFILLER_36_944 VPWR VGND sg13g2_decap_8
XFILLER_35_487 VPWR VGND sg13g2_decap_8
XFILLER_35_498 VPWR VGND sg13g2_decap_8
X_3984_ _0960_ _0943_ _0958_ VPWR VGND sg13g2_xnor2_1
X_5723_ net763 _2488_ _2489_ _0351_ VPWR VGND sg13g2_mux2_1
X_5654_ net476 VPWR _2443_ VGND net586 net1063 sg13g2_o21ai_1
X_4605_ _1512_ _1510_ _1511_ VPWR VGND sg13g2_xnor2_1
Xhold300 mydesign.accum\[33\] VPWR VGND net919 sg13g2_dlygate4sd3_1
Xhold311 mydesign.weights\[3\]\[14\] VPWR VGND net930 sg13g2_dlygate4sd3_1
X_5585_ mydesign.pe_inputs\[6\] net523 mydesign.accum\[2\] _2377_ VPWR VGND sg13g2_nand3_1
XFILLER_11_1024 VPWR VGND sg13g2_decap_4
Xhold322 mydesign.accum\[63\] VPWR VGND net941 sg13g2_dlygate4sd3_1
X_4536_ _1425_ _1446_ _1447_ VPWR VGND sg13g2_nor2b_1
Xhold344 mydesign.accum\[46\] VPWR VGND net963 sg13g2_dlygate4sd3_1
Xhold333 mydesign.pe_weights\[46\] VPWR VGND net952 sg13g2_dlygate4sd3_1
Xhold366 mydesign.weights\[3\]\[12\] VPWR VGND net985 sg13g2_dlygate4sd3_1
Xhold377 mydesign.pe_weights\[54\] VPWR VGND net996 sg13g2_dlygate4sd3_1
Xhold355 mydesign.pe_inputs\[27\] VPWR VGND net974 sg13g2_dlygate4sd3_1
X_4467_ _1389_ VPWR _1391_ VGND _1376_ _1379_ sg13g2_o21ai_1
X_3418_ net516 mydesign.accum\[117\] mydesign.accum\[85\] mydesign.accum\[53\] mydesign.accum\[21\]
+ net508 _0463_ VPWR VGND sg13g2_mux4_1
Xhold388 mydesign.accum\[97\] VPWR VGND net1007 sg13g2_dlygate4sd3_1
X_4398_ _1325_ mydesign.pe_weights\[52\] mydesign.pe_inputs\[43\] VPWR VGND sg13g2_nand2_1
Xhold399 mydesign.accum\[44\] VPWR VGND net1018 sg13g2_dlygate4sd3_1
X_3349_ _0399_ _0401_ _0065_ VPWR VGND sg13g2_nor2_1
X_6137_ net304 VGND VPWR _0363_ mydesign.weights\[0\]\[19\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_46_719 VPWR VGND sg13g2_decap_8
X_6068_ net190 VGND VPWR net641 mydesign.weights\[2\]\[10\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_5019_ _1871_ _1860_ _1862_ VPWR VGND sg13g2_nand2_1
XFILLER_26_410 VPWR VGND sg13g2_fill_1
XFILLER_27_955 VPWR VGND sg13g2_decap_8
XFILLER_42_947 VPWR VGND sg13g2_decap_8
XFILLER_41_402 VPWR VGND sg13g2_decap_4
XFILLER_14_649 VPWR VGND sg13g2_fill_2
XFILLER_6_837 VPWR VGND sg13g2_decap_4
X_6041__294 VPWR VGND net294 sg13g2_tiehi
XFILLER_49_535 VPWR VGND sg13g2_fill_1
XFILLER_45_730 VPWR VGND sg13g2_decap_8
XFILLER_18_988 VPWR VGND sg13g2_decap_8
XFILLER_33_903 VPWR VGND sg13g2_decap_8
XFILLER_44_251 VPWR VGND sg13g2_fill_1
X_5920__317 VPWR VGND net317 sg13g2_tiehi
XFILLER_9_697 VPWR VGND sg13g2_decap_8
X_5370_ _2184_ _2167_ _2185_ VPWR VGND sg13g2_nor2b_1
X_4321_ _1260_ _1240_ _1262_ VPWR VGND sg13g2_xor2_1
X_4252_ mydesign.pe_weights\[58\] net536 mydesign.accum\[82\] _1196_ VPWR VGND sg13g2_nand3_1
XFILLER_4_380 VPWR VGND sg13g2_fill_1
X_3203_ _2634_ VPWR _0009_ VGND _2520_ _2633_ sg13g2_o21ai_1
X_5992__142 VPWR VGND net142 sg13g2_tiehi
X_4183_ _1128_ VPWR _1140_ VGND _1121_ _1129_ sg13g2_o21ai_1
XFILLER_41_1028 VPWR VGND sg13g2_fill_1
X_3134_ VPWR _2575_ net881 VGND sg13g2_inv_1
XFILLER_36_774 VPWR VGND sg13g2_decap_8
XFILLER_23_435 VPWR VGND sg13g2_fill_2
XFILLER_23_457 VPWR VGND sg13g2_fill_2
X_3967_ _0944_ _0941_ _0942_ VPWR VGND sg13g2_xnor2_1
X_5706_ _2480_ VPWR _0343_ VGND net597 _2476_ sg13g2_o21ai_1
X_3898_ _0887_ _0885_ _0886_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_30_clk clknet_3_7__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_5637_ VGND VPWR net586 _2425_ _0328_ _2426_ sg13g2_a21oi_1
X_5568_ net475 VPWR _2362_ VGND net749 _2361_ sg13g2_o21ai_1
Xhold130 mydesign.accum\[0\] VPWR VGND net749 sg13g2_dlygate4sd3_1
X_4519_ _1413_ _1429_ _1431_ VPWR VGND sg13g2_nor2_1
Xhold152 mydesign.weights\[1\]\[12\] VPWR VGND net771 sg13g2_dlygate4sd3_1
Xhold141 mydesign.inputs\[0\]\[25\] VPWR VGND net760 sg13g2_dlygate4sd3_1
Xhold174 mydesign.inputs\[1\]\[22\] VPWR VGND net793 sg13g2_dlygate4sd3_1
Xhold163 mydesign.inputs\[1\]\[17\] VPWR VGND net782 sg13g2_dlygate4sd3_1
Xhold185 mydesign.accum\[91\] VPWR VGND net804 sg13g2_dlygate4sd3_1
X_5499_ _2301_ _2299_ _2300_ VPWR VGND sg13g2_nand2_1
Xfanout610 net611 net610 VPWR VGND sg13g2_buf_8
Xfanout632 net639 net632 VPWR VGND sg13g2_buf_8
Xfanout621 net640 net621 VPWR VGND sg13g2_buf_8
Xhold196 mydesign.pe_weights\[44\] VPWR VGND net815 sg13g2_dlygate4sd3_1
X_5971__215 VPWR VGND net215 sg13g2_tiehi
XFILLER_37_44 VPWR VGND sg13g2_decap_4
XFILLER_41_221 VPWR VGND sg13g2_decap_8
XFILLER_15_958 VPWR VGND sg13g2_decap_8
XFILLER_30_906 VPWR VGND sg13g2_decap_8
XFILLER_23_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_21_clk clknet_3_3__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_6_645 VPWR VGND sg13g2_decap_8
XFILLER_49_310 VPWR VGND sg13g2_decap_4
XFILLER_49_365 VPWR VGND sg13g2_fill_1
XFILLER_49_354 VPWR VGND sg13g2_decap_4
X_4870_ VGND VPWR _1727_ _1730_ _1746_ _1745_ sg13g2_a21oi_1
X_3821_ mydesign.pe_inputs\[56\] _0783_ net688 _0814_ VPWR VGND sg13g2_nand3_1
XFILLER_21_939 VPWR VGND sg13g2_decap_8
XFILLER_14_991 VPWR VGND sg13g2_decap_8
XFILLER_32_276 VPWR VGND sg13g2_fill_2
XFILLER_32_287 VPWR VGND sg13g2_fill_1
X_3752_ _0756_ _0758_ _0742_ _0760_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_12_clk clknet_3_2__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_3683_ _0691_ _0692_ _0693_ _0694_ VPWR VGND sg13g2_or3_1
X_5422_ _2220_ _2223_ _2233_ _2234_ VPWR VGND sg13g2_or3_1
X_5353_ _2159_ VPWR _2168_ VGND _2152_ _2160_ sg13g2_o21ai_1
X_4304_ _1225_ _1227_ _1245_ _1246_ VPWR VGND sg13g2_nor3_1
X_6055__238 VPWR VGND net238 sg13g2_tiehi
X_5284_ mydesign.pe_weights\[31\] _2020_ mydesign.accum\[30\] _2112_ VPWR VGND sg13g2_nand3_1
X_4235_ VGND VPWR _2564_ net448 _0171_ _1181_ sg13g2_a21oi_1
X_4166_ mydesign.pe_weights\[63\] _1051_ _1124_ VPWR VGND sg13g2_and2_1
X_3117_ VPWR _2558_ net971 VGND sg13g2_inv_1
X_4097_ net624 VPWR _1063_ VGND net815 net436 sg13g2_o21ai_1
XFILLER_24_700 VPWR VGND sg13g2_decap_8
XFILLER_24_711 VPWR VGND sg13g2_fill_2
XFILLER_24_755 VPWR VGND sg13g2_fill_2
XFILLER_36_582 VPWR VGND sg13g2_decap_4
XFILLER_12_906 VPWR VGND sg13g2_fill_2
XFILLER_12_928 VPWR VGND sg13g2_decap_8
XFILLER_23_243 VPWR VGND sg13g2_fill_2
X_4999_ net477 VPWR _1853_ VGND net585 net1018 sg13g2_o21ai_1
XFILLER_20_961 VPWR VGND sg13g2_decap_8
XFILLER_23_68 VPWR VGND sg13g2_decap_8
XFILLER_48_32 VPWR VGND sg13g2_fill_1
XFILLER_48_21 VPWR VGND sg13g2_decap_8
Xfanout440 net441 net440 VPWR VGND sg13g2_buf_8
XFILLER_47_803 VPWR VGND sg13g2_decap_8
Xfanout484 net485 net484 VPWR VGND sg13g2_buf_8
Xfanout473 net474 net473 VPWR VGND sg13g2_buf_8
Xfanout462 _2661_ net462 VPWR VGND sg13g2_buf_8
XFILLER_24_1023 VPWR VGND sg13g2_decap_4
Xfanout451 net452 net451 VPWR VGND sg13g2_buf_8
XFILLER_48_87 VPWR VGND sg13g2_fill_2
Xfanout495 net496 net495 VPWR VGND sg13g2_buf_8
XFILLER_46_368 VPWR VGND sg13g2_decap_8
XFILLER_27_571 VPWR VGND sg13g2_decap_8
XFILLER_15_733 VPWR VGND sg13g2_decap_8
XFILLER_30_725 VPWR VGND sg13g2_decap_4
XFILLER_11_961 VPWR VGND sg13g2_decap_8
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_140 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_1_clk clknet_3_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
X_4020_ _0993_ _0990_ _0994_ VPWR VGND sg13g2_xor2_1
XFILLER_49_184 VPWR VGND sg13g2_fill_1
XFILLER_37_357 VPWR VGND sg13g2_decap_4
XFILLER_46_880 VPWR VGND sg13g2_decap_8
X_5971_ net215 VGND VPWR _0197_ mydesign.inputs\[3\]\[13\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_4922_ VGND VPWR _2535_ net445 _0257_ _1782_ sg13g2_a21oi_1
X_4853_ VGND VPWR _1730_ _1729_ _1726_ sg13g2_or2_1
XFILLER_21_725 VPWR VGND sg13g2_fill_1
XFILLER_33_585 VPWR VGND sg13g2_fill_2
X_3804_ net550 mydesign.weights\[2\]\[11\] _0799_ VPWR VGND sg13g2_nor2_1
XFILLER_20_235 VPWR VGND sg13g2_fill_1
XFILLER_21_769 VPWR VGND sg13g2_fill_1
X_4784_ mydesign.pe_weights\[40\] net529 net745 _1665_ VPWR VGND _1663_ sg13g2_nand4_1
X_3735_ _0744_ _0721_ _0741_ VPWR VGND sg13g2_xnor2_1
X_5405_ _2218_ _2216_ _2217_ VPWR VGND sg13g2_nand2_1
X_3666_ _0674_ _0675_ _0677_ _0678_ VPWR VGND sg13g2_nor3_1
X_3597_ _0606_ _0620_ _0621_ VPWR VGND sg13g2_nor2_1
XFILLER_0_629 VPWR VGND sg13g2_decap_8
X_5336_ _2152_ mydesign.pe_inputs\[14\] mydesign.pe_weights\[24\] VPWR VGND sg13g2_nand2_1
X_5267_ _2096_ mydesign.pe_weights\[30\] _2020_ VPWR VGND sg13g2_nand2_1
X_4218_ net471 VPWR _1173_ VGND net569 net948 sg13g2_o21ai_1
X_5864__45 VPWR VGND net45 sg13g2_tiehi
X_5198_ _2031_ mydesign.accum\[24\] _2022_ _2030_ VPWR VGND sg13g2_and3_2
X_4149_ _1100_ _1106_ _1107_ _1108_ VPWR VGND sg13g2_or3_1
XFILLER_44_806 VPWR VGND sg13g2_decap_8
XFILLER_28_368 VPWR VGND sg13g2_decap_4
XFILLER_34_56 VPWR VGND sg13g2_decap_8
Xheichips25_template_405 VPWR VGND uio_oe[6] sg13g2_tiehi
Xclkload0 clknet_3_1__leaf_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_1_2 VPWR VGND sg13g2_fill_1
XFILLER_47_600 VPWR VGND sg13g2_decap_8
XFILLER_35_806 VPWR VGND sg13g2_decap_8
XFILLER_47_677 VPWR VGND sg13g2_decap_8
XFILLER_46_198 VPWR VGND sg13g2_fill_1
XFILLER_43_872 VPWR VGND sg13g2_decap_8
XFILLER_15_574 VPWR VGND sg13g2_decap_8
XFILLER_15_585 VPWR VGND sg13g2_fill_1
X_5884__381 VPWR VGND net381 sg13g2_tiehi
X_3520_ _0548_ _0530_ _0546_ VPWR VGND sg13g2_xnor2_1
X_3451_ VGND VPWR net607 _0493_ _0491_ net606 sg13g2_a21oi_2
X_3382_ net511 mydesign.accum\[122\] mydesign.accum\[90\] mydesign.accum\[58\] mydesign.accum\[26\]
+ net505 _0430_ VPWR VGND sg13g2_mux4_1
X_5121_ _1961_ _1962_ _0276_ VPWR VGND sg13g2_nor2_1
XFILLER_38_611 VPWR VGND sg13g2_fill_2
X_5052_ VGND VPWR mydesign.pe_weights\[33\] net526 _1897_ mydesign.accum\[33\] sg13g2_a21oi_1
X_4003_ _0975_ _0976_ _0953_ _0978_ VPWR VGND sg13g2_nand3_1
XFILLER_37_143 VPWR VGND sg13g2_fill_1
XFILLER_19_880 VPWR VGND sg13g2_fill_2
XFILLER_19_891 VPWR VGND sg13g2_fill_2
X_5954_ net249 VGND VPWR _0180_ mydesign.pe_inputs\[36\] clknet_leaf_40_clk sg13g2_dfrbpq_2
X_5885_ net379 VGND VPWR _0111_ mydesign.accum\[119\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_4905_ _1773_ net3 _1768_ VPWR VGND sg13g2_nand2_2
XFILLER_21_544 VPWR VGND sg13g2_fill_2
X_4836_ _1713_ _1704_ _1714_ VPWR VGND sg13g2_xor2_1
X_4767_ VGND VPWR _2544_ net451 _0232_ _1652_ sg13g2_a21oi_1
X_4698_ VGND VPWR net560 _1591_ _0223_ _1592_ sg13g2_a21oi_1
X_3718_ _0728_ _0725_ _0726_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_47 VPWR VGND sg13g2_fill_2
X_3649_ net463 _0662_ _0104_ VPWR VGND sg13g2_nor2_1
X_5319_ VGND VPWR _2526_ net449 _0298_ _2138_ sg13g2_a21oi_1
XFILLER_49_909 VPWR VGND sg13g2_decap_8
XFILLER_0_459 VPWR VGND sg13g2_fill_2
Xhold12 mydesign.inputs\[2\]\[14\] VPWR VGND net418 sg13g2_dlygate4sd3_1
Xhold23 mydesign.inputs\[2\]\[11\] VPWR VGND net642 sg13g2_dlygate4sd3_1
Xhold45 mydesign.accum\[40\] VPWR VGND net664 sg13g2_dlygate4sd3_1
Xhold56 mydesign.weights\[2\]\[17\] VPWR VGND net675 sg13g2_dlygate4sd3_1
Xhold34 _0079_ VPWR VGND net653 sg13g2_dlygate4sd3_1
Xhold89 _0115_ VPWR VGND net708 sg13g2_dlygate4sd3_1
Xhold78 mydesign.inputs\[3\]\[5\] VPWR VGND net697 sg13g2_dlygate4sd3_1
Xhold67 mydesign.accum\[56\] VPWR VGND net686 sg13g2_dlygate4sd3_1
XFILLER_44_603 VPWR VGND sg13g2_fill_1
XFILLER_17_806 VPWR VGND sg13g2_fill_1
XFILLER_17_839 VPWR VGND sg13g2_decap_8
X_6014__34 VPWR VGND net34 sg13g2_tiehi
XFILLER_24_360 VPWR VGND sg13g2_fill_2
XFILLER_25_883 VPWR VGND sg13g2_fill_2
X_6148__272 VPWR VGND net272 sg13g2_tiehi
XFILLER_12_533 VPWR VGND sg13g2_fill_2
XFILLER_40_875 VPWR VGND sg13g2_decap_8
XFILLER_4_721 VPWR VGND sg13g2_fill_1
XFILLER_0_971 VPWR VGND sg13g2_decap_8
XFILLER_48_986 VPWR VGND sg13g2_decap_8
XFILLER_34_124 VPWR VGND sg13g2_fill_2
XFILLER_43_680 VPWR VGND sg13g2_decap_8
XFILLER_37_1022 VPWR VGND sg13g2_decap_8
XFILLER_34_168 VPWR VGND sg13g2_fill_2
XFILLER_42_190 VPWR VGND sg13g2_fill_1
X_5670_ VGND VPWR _2444_ _2450_ _2457_ _2453_ sg13g2_a21oi_1
X_4621_ net460 VPWR _1526_ VGND net557 mydesign.inputs\[2\]\[9\] sg13g2_o21ai_1
XFILLER_30_396 VPWR VGND sg13g2_decap_4
X_4552_ net537 mydesign.pe_inputs\[37\] mydesign.accum\[68\] _1462_ VPWR VGND sg13g2_nand3_1
X_4483_ _1404_ net644 _1402_ VPWR VGND sg13g2_nand2_1
X_3503_ _0532_ _0530_ _0531_ VPWR VGND sg13g2_nand2_1
X_3434_ VPWR VGND net458 _0477_ _0472_ _0412_ _0478_ _0471_ sg13g2_a221oi_1
X_3365_ VGND VPWR net456 _0408_ _0415_ _2698_ sg13g2_a21oi_1
X_3296_ _2668_ net786 _2690_ _0046_ VPWR VGND sg13g2_mux2_1
X_5104_ mydesign.pe_inputs\[22\] net530 mydesign.accum\[36\] _1946_ VPWR VGND sg13g2_a21o_1
X_6084_ net36 VGND VPWR net833 mydesign.pe_inputs\[6\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_39_942 VPWR VGND sg13g2_decap_8
X_5035_ _1872_ net980 _1886_ VPWR VGND sg13g2_xor2_1
XFILLER_38_496 VPWR VGND sg13g2_decap_4
X_5937_ net283 VGND VPWR _0163_ mydesign.accum\[95\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_5868_ net37 VGND VPWR _0094_ mydesign.accum\[126\] clknet_leaf_16_clk sg13g2_dfrbpq_2
XFILLER_21_352 VPWR VGND sg13g2_decap_8
X_4819_ _1697_ _1685_ _1698_ VPWR VGND sg13g2_xor2_1
X_5799_ net151 VGND VPWR _0025_ mydesign.inputs\[1\]\[12\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_5_529 VPWR VGND sg13g2_decap_8
Xoutput13 net13 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_735 VPWR VGND sg13g2_fill_2
XFILLER_49_706 VPWR VGND sg13g2_decap_8
XFILLER_45_912 VPWR VGND sg13g2_decap_8
XFILLER_17_614 VPWR VGND sg13g2_fill_1
XFILLER_45_989 VPWR VGND sg13g2_decap_8
XFILLER_17_658 VPWR VGND sg13g2_decap_8
XFILLER_40_661 VPWR VGND sg13g2_decap_8
XFILLER_9_824 VPWR VGND sg13g2_decap_4
XFILLER_12_341 VPWR VGND sg13g2_fill_2
XFILLER_8_334 VPWR VGND sg13g2_fill_1
XFILLER_8_323 VPWR VGND sg13g2_decap_8
XFILLER_9_879 VPWR VGND sg13g2_fill_1
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_39_216 VPWR VGND sg13g2_fill_1
X_3150_ _2591_ net610 VPWR VGND sg13g2_inv_8
X_3081_ VPWR _2522_ net832 VGND sg13g2_inv_1
XFILLER_11_4 VPWR VGND sg13g2_decap_8
XFILLER_48_783 VPWR VGND sg13g2_decap_8
XFILLER_47_282 VPWR VGND sg13g2_fill_1
XFILLER_36_923 VPWR VGND sg13g2_decap_8
XFILLER_35_444 VPWR VGND sg13g2_fill_1
XFILLER_23_639 VPWR VGND sg13g2_fill_2
X_3983_ _0959_ _0943_ _0958_ VPWR VGND sg13g2_nand2_1
X_5722_ net761 _2487_ _2489_ _0350_ VPWR VGND sg13g2_mux2_1
X_5653_ _2442_ _2427_ _2440_ VPWR VGND sg13g2_xnor2_1
X_5584_ _2376_ mydesign.accum\[2\] mydesign.pe_inputs\[6\] net523 VPWR VGND sg13g2_and3_1
X_4604_ _1511_ net843 _1497_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_1003 VPWR VGND sg13g2_decap_8
XFILLER_8_890 VPWR VGND sg13g2_fill_2
Xhold301 _0273_ VPWR VGND net920 sg13g2_dlygate4sd3_1
X_4535_ _1445_ _1442_ _1446_ VPWR VGND sg13g2_xor2_1
Xhold312 _2508_ VPWR VGND net931 sg13g2_dlygate4sd3_1
Xhold323 mydesign.accum\[109\] VPWR VGND net942 sg13g2_dlygate4sd3_1
Xhold334 _0218_ VPWR VGND net953 sg13g2_dlygate4sd3_1
Xhold378 mydesign.accum\[92\] VPWR VGND net997 sg13g2_dlygate4sd3_1
Xhold345 mydesign.accum\[90\] VPWR VGND net964 sg13g2_dlygate4sd3_1
Xhold356 _0255_ VPWR VGND net975 sg13g2_dlygate4sd3_1
Xhold367 _2506_ VPWR VGND net986 sg13g2_dlygate4sd3_1
X_4466_ _1376_ _1379_ _1389_ _1390_ VPWR VGND sg13g2_or3_1
Xhold389 _0141_ VPWR VGND net1008 sg13g2_dlygate4sd3_1
X_4397_ _1315_ VPWR _1324_ VGND _1308_ _1316_ sg13g2_o21ai_1
X_3417_ net430 VPWR _0462_ VGND _0460_ _0461_ sg13g2_o21ai_1
X_3348_ _0401_ net619 _0400_ VPWR VGND sg13g2_nand2_1
X_6136_ net312 VGND VPWR _0362_ mydesign.weights\[0\]\[18\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3279_ _2683_ mydesign.load_counter\[0\] VPWR VGND mydesign.load_counter\[1\] sg13g2_nand2b_2
X_6067_ net192 VGND VPWR net661 mydesign.weights\[2\]\[9\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_39_783 VPWR VGND sg13g2_fill_1
X_5018_ net463 _1870_ _0265_ VPWR VGND sg13g2_nor2_1
XFILLER_27_934 VPWR VGND sg13g2_decap_8
XFILLER_42_926 VPWR VGND sg13g2_decap_8
XFILLER_14_606 VPWR VGND sg13g2_decap_8
XFILLER_14_639 VPWR VGND sg13g2_fill_2
XFILLER_26_477 VPWR VGND sg13g2_fill_2
XFILLER_26_499 VPWR VGND sg13g2_decap_8
XFILLER_9_109 VPWR VGND sg13g2_fill_2
XFILLER_42_45 VPWR VGND sg13g2_fill_1
XFILLER_22_672 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_fill_2
XFILLER_49_547 VPWR VGND sg13g2_decap_8
XFILLER_18_967 VPWR VGND sg13g2_decap_8
XFILLER_45_786 VPWR VGND sg13g2_decap_8
XFILLER_33_959 VPWR VGND sg13g2_decap_8
XFILLER_32_458 VPWR VGND sg13g2_fill_1
XFILLER_8_131 VPWR VGND sg13g2_decap_8
X_4320_ _1240_ _1260_ _1261_ VPWR VGND sg13g2_nor2b_1
X_4251_ _1195_ mydesign.pe_weights\[57\] mydesign.pe_inputs\[45\] VPWR VGND sg13g2_nand2_1
X_3202_ net617 _2633_ net677 _2634_ VPWR VGND sg13g2_nand3_1
X_4182_ VGND VPWR _1134_ _1136_ _1139_ _1133_ sg13g2_a21oi_1
XFILLER_41_1007 VPWR VGND sg13g2_decap_8
X_3133_ VPWR _2574_ net804 VGND sg13g2_inv_1
XFILLER_36_720 VPWR VGND sg13g2_decap_8
XFILLER_24_904 VPWR VGND sg13g2_fill_2
X_3966_ _0941_ _0942_ _0943_ VPWR VGND sg13g2_nor2b_1
X_5705_ net731 _2476_ net613 _2480_ VPWR VGND sg13g2_nand3_1
XFILLER_32_992 VPWR VGND sg13g2_decap_8
X_5636_ net476 VPWR _2426_ VGND net586 net1068 sg13g2_o21ai_1
X_3897_ _0864_ _0866_ _0884_ _0886_ VPWR VGND sg13g2_or3_1
X_5567_ _2361_ net587 mydesign.pe_inputs\[4\] mydesign.pe_weights\[16\] VPWR VGND
+ sg13g2_and3_1
Xhold153 mydesign.inputs\[0\]\[14\] VPWR VGND net772 sg13g2_dlygate4sd3_1
Xhold120 mydesign.accum\[80\] VPWR VGND net739 sg13g2_dlygate4sd3_1
Xhold131 _0324_ VPWR VGND net750 sg13g2_dlygate4sd3_1
XFILLER_2_318 VPWR VGND sg13g2_decap_4
X_4518_ _1430_ _1413_ _1429_ VPWR VGND sg13g2_nand2_1
X_5498_ net525 mydesign.pe_inputs\[10\] mydesign.accum\[12\] _2300_ VPWR VGND sg13g2_a21o_1
Xhold142 mydesign.weights\[1\]\[14\] VPWR VGND net761 sg13g2_dlygate4sd3_1
Xhold186 mydesign.weights\[2\]\[12\] VPWR VGND net805 sg13g2_dlygate4sd3_1
X_4449_ _1374_ _1372_ _1373_ VPWR VGND sg13g2_nand2_1
Xhold164 mydesign.inputs\[0\]\[20\] VPWR VGND net783 sg13g2_dlygate4sd3_1
Xhold175 mydesign.inputs\[1\]\[8\] VPWR VGND net794 sg13g2_dlygate4sd3_1
Xhold197 mydesign.pe_weights\[35\] VPWR VGND net816 sg13g2_dlygate4sd3_1
Xfanout633 net636 net633 VPWR VGND sg13g2_buf_8
Xfanout611 ui_in[4] net611 VPWR VGND sg13g2_buf_8
Xfanout622 net623 net622 VPWR VGND sg13g2_buf_8
Xfanout600 _2629_ net600 VPWR VGND sg13g2_buf_8
X_5819__123 VPWR VGND net123 sg13g2_tiehi
X_6119_ net84 VGND VPWR _0345_ mydesign.weights\[1\]\[9\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_27_731 VPWR VGND sg13g2_fill_2
XFILLER_42_701 VPWR VGND sg13g2_fill_1
XFILLER_15_937 VPWR VGND sg13g2_decap_8
XFILLER_27_764 VPWR VGND sg13g2_decap_8
XFILLER_27_797 VPWR VGND sg13g2_fill_2
XFILLER_42_745 VPWR VGND sg13g2_decap_8
XFILLER_18_1009 VPWR VGND sg13g2_decap_8
XFILLER_26_296 VPWR VGND sg13g2_fill_2
XFILLER_42_767 VPWR VGND sg13g2_decap_8
X_5826__116 VPWR VGND net116 sg13g2_tiehi
XFILLER_10_653 VPWR VGND sg13g2_decap_4
XFILLER_2_896 VPWR VGND sg13g2_decap_8
XFILLER_1_373 VPWR VGND sg13g2_fill_1
XFILLER_37_528 VPWR VGND sg13g2_fill_1
XFILLER_18_731 VPWR VGND sg13g2_fill_1
XFILLER_45_561 VPWR VGND sg13g2_decap_8
X_3820_ _0811_ _0810_ _0813_ VPWR VGND sg13g2_xor2_1
XFILLER_33_778 VPWR VGND sg13g2_fill_2
X_3751_ _0758_ _0742_ _0756_ _0759_ VPWR VGND sg13g2_a21o_1
XFILLER_14_970 VPWR VGND sg13g2_decap_8
X_3682_ VGND VPWR net540 _0658_ _0693_ mydesign.accum\[115\] sg13g2_a21oi_1
X_5421_ _2233_ _2231_ _2232_ VPWR VGND sg13g2_xnor2_1
X_5352_ _2163_ VPWR _2167_ VGND _2149_ _2164_ sg13g2_o21ai_1
X_4303_ _1243_ _1242_ _1245_ VPWR VGND sg13g2_xor2_1
X_5283_ VGND VPWR mydesign.pe_weights\[31\] _2020_ _2111_ mydesign.accum\[30\] sg13g2_a21oi_1
X_4234_ net631 VPWR _1181_ VGND net533 net448 sg13g2_o21ai_1
X_4165_ _1123_ mydesign.pe_weights\[62\] _1056_ VPWR VGND sg13g2_nand2_1
X_3116_ VPWR _2557_ net996 VGND sg13g2_inv_1
X_4096_ VGND VPWR _2568_ net488 _0151_ _1062_ sg13g2_a21oi_1
XFILLER_24_778 VPWR VGND sg13g2_fill_1
XFILLER_17_1020 VPWR VGND sg13g2_decap_8
X_4998_ VGND VPWR _1850_ _1851_ _1852_ net501 sg13g2_a21oi_1
X_3949_ _0928_ mydesign.weights\[3\]\[11\] net548 VPWR VGND sg13g2_nand2b_1
XFILLER_20_940 VPWR VGND sg13g2_decap_8
X_5619_ _2397_ VPWR _2409_ VGND _2389_ _2398_ sg13g2_o21ai_1
Xfanout441 net453 net441 VPWR VGND sg13g2_buf_8
Xfanout430 net431 net430 VPWR VGND sg13g2_buf_8
XFILLER_24_1002 VPWR VGND sg13g2_decap_8
Xfanout474 net478 net474 VPWR VGND sg13g2_buf_8
Xfanout463 _2661_ net463 VPWR VGND sg13g2_buf_8
Xfanout452 net453 net452 VPWR VGND sg13g2_buf_8
XFILLER_46_314 VPWR VGND sg13g2_fill_1
Xfanout496 _2595_ net496 VPWR VGND sg13g2_buf_8
Xfanout485 _2602_ net485 VPWR VGND sg13g2_buf_8
XFILLER_47_859 VPWR VGND sg13g2_decap_8
XFILLER_42_553 VPWR VGND sg13g2_fill_2
XFILLER_14_288 VPWR VGND sg13g2_fill_1
XFILLER_30_715 VPWR VGND sg13g2_fill_1
XFILLER_11_940 VPWR VGND sg13g2_decap_8
XFILLER_31_1006 VPWR VGND sg13g2_decap_8
XFILLER_10_472 VPWR VGND sg13g2_fill_1
XFILLER_7_988 VPWR VGND sg13g2_decap_8
XFILLER_43_7 VPWR VGND sg13g2_fill_1
XFILLER_49_163 VPWR VGND sg13g2_decap_8
XFILLER_49_196 VPWR VGND sg13g2_decap_4
XFILLER_38_859 VPWR VGND sg13g2_fill_2
X_5970_ net217 VGND VPWR _0196_ mydesign.inputs\[3\]\[12\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_6089__368 VPWR VGND net368 sg13g2_tiehi
XFILLER_45_380 VPWR VGND sg13g2_fill_1
X_4921_ net635 VPWR _1782_ VGND mydesign.pe_weights\[21\] net445 sg13g2_o21ai_1
X_4852_ _1729_ _1727_ _1728_ VPWR VGND sg13g2_nand2_1
X_3803_ mydesign.weights\[2\]\[7\] net551 _0798_ VPWR VGND sg13g2_nor2b_1
X_4783_ mydesign.pe_weights\[40\] net529 net745 _1664_ VPWR VGND sg13g2_nand3_1
X_3734_ _0721_ _0741_ _0743_ VPWR VGND sg13g2_nor2_1
X_3665_ _0677_ mydesign.pe_inputs\[61\] _0648_ VPWR VGND sg13g2_nand2_1
X_5404_ _2195_ VPWR _2217_ VGND _2188_ _2196_ sg13g2_o21ai_1
XFILLER_47_1013 VPWR VGND sg13g2_decap_8
X_3596_ _0620_ _0615_ _0619_ VPWR VGND sg13g2_xnor2_1
X_5335_ VGND VPWR net591 _2150_ _0301_ _2151_ sg13g2_a21oi_1
X_5266_ _2085_ VPWR _2095_ VGND _2078_ _2086_ sg13g2_o21ai_1
X_4217_ _1172_ _1168_ _1171_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_25 VPWR VGND sg13g2_fill_1
X_5197_ _2028_ _2027_ _2030_ VPWR VGND sg13g2_xor2_1
X_4148_ VGND VPWR _1104_ _1105_ _1107_ _1081_ sg13g2_a21oi_1
X_5816__126 VPWR VGND net126 sg13g2_tiehi
XFILLER_37_870 VPWR VGND sg13g2_fill_2
X_4079_ mydesign.inputs\[1\]\[9\] net460 net498 _1048_ VPWR VGND sg13g2_nand3_1
XFILLER_24_553 VPWR VGND sg13g2_decap_4
XFILLER_11_203 VPWR VGND sg13g2_fill_2
XFILLER_11_236 VPWR VGND sg13g2_fill_2
Xheichips25_template_406 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_11_258 VPWR VGND sg13g2_fill_1
Xclkload1 clknet_3_2__leaf_clk clkload1/X VPWR VGND sg13g2_buf_8
X_5823__119 VPWR VGND net119 sg13g2_tiehi
XFILLER_4_925 VPWR VGND sg13g2_fill_1
XFILLER_4_969 VPWR VGND sg13g2_decap_8
XFILLER_47_656 VPWR VGND sg13g2_decap_8
XFILLER_43_851 VPWR VGND sg13g2_decap_8
XFILLER_15_531 VPWR VGND sg13g2_decap_4
XFILLER_15_553 VPWR VGND sg13g2_fill_2
XFILLER_30_501 VPWR VGND sg13g2_fill_1
X_3450_ _0492_ net606 _0491_ VPWR VGND sg13g2_nand2_2
X_3381_ net513 mydesign.accum\[106\] mydesign.accum\[74\] mydesign.accum\[42\] mydesign.accum\[10\]
+ net506 _0429_ VPWR VGND sg13g2_mux4_1
X_5120_ net475 VPWR _1962_ VGND net584 net1002 sg13g2_o21ai_1
X_5051_ _1896_ mydesign.accum\[33\] mydesign.pe_weights\[33\] net526 VPWR VGND sg13g2_and3_2
X_4002_ _0975_ _0976_ _0977_ VPWR VGND sg13g2_and2_1
XFILLER_37_155 VPWR VGND sg13g2_fill_2
X_5953_ net251 VGND VPWR _0179_ mydesign.accum\[87\] clknet_leaf_25_clk sg13g2_dfrbpq_2
XFILLER_40_309 VPWR VGND sg13g2_fill_2
X_5884_ net381 VGND VPWR _0110_ mydesign.accum\[118\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4904_ VGND VPWR _1767_ _1771_ _0249_ net859 sg13g2_a21oi_1
X_4835_ _1713_ _1705_ _1711_ VPWR VGND sg13g2_xnor2_1
XFILLER_14_1012 VPWR VGND sg13g2_decap_8
X_4766_ net637 VPWR _1652_ VGND mydesign.pe_weights\[24\] net451 sg13g2_o21ai_1
X_3717_ _0725_ _0726_ _0727_ VPWR VGND sg13g2_nor2_1
X_4697_ net467 VPWR _1592_ VGND net560 net990 sg13g2_o21ai_1
X_3648_ _0661_ net991 _0662_ VPWR VGND sg13g2_xor2_1
X_3579_ _0602_ _0600_ _0604_ VPWR VGND sg13g2_xor2_1
X_5318_ net638 VPWR _2138_ VGND net832 net449 sg13g2_o21ai_1
XFILLER_0_438 VPWR VGND sg13g2_decap_8
Xhold13 _0078_ VPWR VGND net419 sg13g2_dlygate4sd3_1
X_5937__283 VPWR VGND net283 sg13g2_tiehi
Xhold35 mydesign.inputs\[3\]\[4\] VPWR VGND net654 sg13g2_dlygate4sd3_1
Xhold46 _0260_ VPWR VGND net665 sg13g2_dlygate4sd3_1
Xhold24 _0016_ VPWR VGND net643 sg13g2_dlygate4sd3_1
X_5249_ _2079_ _2057_ _2059_ VPWR VGND sg13g2_nand2_1
Xhold79 mydesign.weights\[0\]\[18\] VPWR VGND net698 sg13g2_dlygate4sd3_1
Xhold57 _0010_ VPWR VGND net676 sg13g2_dlygate4sd3_1
XFILLER_21_1016 VPWR VGND sg13g2_decap_8
XFILLER_21_1027 VPWR VGND sg13g2_fill_2
Xhold68 _0220_ VPWR VGND net687 sg13g2_dlygate4sd3_1
XFILLER_16_306 VPWR VGND sg13g2_fill_1
XFILLER_28_133 VPWR VGND sg13g2_fill_2
XFILLER_16_339 VPWR VGND sg13g2_decap_4
XFILLER_44_659 VPWR VGND sg13g2_decap_8
XFILLER_40_821 VPWR VGND sg13g2_fill_1
XFILLER_12_512 VPWR VGND sg13g2_decap_8
XFILLER_8_527 VPWR VGND sg13g2_decap_8
X_6044__282 VPWR VGND net282 sg13g2_tiehi
XFILLER_3_265 VPWR VGND sg13g2_decap_4
XFILLER_3_298 VPWR VGND sg13g2_fill_2
XFILLER_0_950 VPWR VGND sg13g2_decap_8
XFILLER_48_965 VPWR VGND sg13g2_decap_8
XFILLER_37_1001 VPWR VGND sg13g2_decap_8
XFILLER_35_659 VPWR VGND sg13g2_fill_1
X_4620_ net498 mydesign.inputs\[2\]\[5\] _1525_ VPWR VGND sg13g2_nor2_1
XFILLER_31_887 VPWR VGND sg13g2_decap_8
X_4551_ _1461_ mydesign.pe_weights\[50\] mydesign.pe_inputs\[38\] VPWR VGND sg13g2_nand2_1
XFILLER_7_571 VPWR VGND sg13g2_decap_8
X_4482_ _1403_ VPWR _0196_ VGND net603 _1401_ sg13g2_o21ai_1
X_3502_ _0520_ net455 mydesign.accum\[121\] _0531_ VPWR VGND sg13g2_a21o_1
X_3433_ VGND VPWR net509 _0475_ _0477_ _0476_ sg13g2_a21oi_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
XFILLER_44_1016 VPWR VGND sg13g2_decap_8
X_5103_ net530 mydesign.pe_inputs\[22\] mydesign.accum\[36\] _1945_ VPWR VGND sg13g2_nand3_1
X_6134__328 VPWR VGND net328 sg13g2_tiehi
X_3364_ VGND VPWR net507 _0411_ _0414_ _0413_ sg13g2_a21oi_1
XFILLER_39_921 VPWR VGND sg13g2_decap_8
X_6083_ net44 VGND VPWR net935 mydesign.pe_inputs\[5\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3295_ _2667_ net765 _2690_ _0045_ VPWR VGND sg13g2_mux2_1
X_5034_ VGND VPWR _1860_ _1877_ _1885_ _1876_ sg13g2_a21oi_1
X_5813__129 VPWR VGND net129 sg13g2_tiehi
XFILLER_39_998 VPWR VGND sg13g2_decap_8
XFILLER_25_125 VPWR VGND sg13g2_fill_2
X_5936_ net285 VGND VPWR _0162_ mydesign.accum\[94\] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_22_810 VPWR VGND sg13g2_decap_4
XFILLER_34_692 VPWR VGND sg13g2_fill_2
X_5867_ net39 VGND VPWR _0093_ mydesign.accum\[125\] clknet_leaf_16_clk sg13g2_dfrbpq_2
XFILLER_21_331 VPWR VGND sg13g2_fill_1
XFILLER_22_865 VPWR VGND sg13g2_fill_1
X_5798_ net152 VGND VPWR _0024_ mydesign.inputs\[1\]\[11\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_4818_ _1697_ _1673_ _1695_ VPWR VGND sg13g2_xnor2_1
X_4749_ net470 VPWR _1641_ VGND net567 net884 sg13g2_o21ai_1
XFILLER_5_519 VPWR VGND sg13g2_decap_4
Xoutput14 net14 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_213 VPWR VGND sg13g2_decap_4
XFILLER_5_1021 VPWR VGND sg13g2_decap_8
XFILLER_45_968 VPWR VGND sg13g2_decap_8
XFILLER_4_530 VPWR VGND sg13g2_fill_2
X_3080_ VPWR _2521_ net520 VGND sg13g2_inv_1
XFILLER_48_762 VPWR VGND sg13g2_decap_8
XFILLER_36_902 VPWR VGND sg13g2_decap_8
XFILLER_35_423 VPWR VGND sg13g2_decap_4
XFILLER_36_979 VPWR VGND sg13g2_decap_8
X_3982_ _0958_ _0949_ _0956_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_607 VPWR VGND sg13g2_fill_2
XFILLER_23_618 VPWR VGND sg13g2_decap_8
XFILLER_22_139 VPWR VGND sg13g2_fill_2
X_5721_ net764 _2486_ _2489_ _0349_ VPWR VGND sg13g2_mux2_1
X_5652_ _2441_ _2427_ _2440_ VPWR VGND sg13g2_nand2_1
XFILLER_31_695 VPWR VGND sg13g2_decap_8
X_5583_ _2375_ mydesign.pe_inputs\[5\] mydesign.pe_weights\[17\] VPWR VGND sg13g2_nand2_1
X_4603_ VGND VPWR _1486_ _1501_ _1510_ _1500_ sg13g2_a21oi_1
X_4534_ _1445_ _1443_ _1444_ VPWR VGND sg13g2_nand2_1
Xhold302 mydesign.accum\[42\] VPWR VGND net921 sg13g2_dlygate4sd3_1
Xhold313 _0366_ VPWR VGND net932 sg13g2_dlygate4sd3_1
Xhold324 mydesign.pe_weights\[36\] VPWR VGND net943 sg13g2_dlygate4sd3_1
X_6058__226 VPWR VGND net226 sg13g2_tiehi
Xhold335 mydesign.accum\[25\] VPWR VGND net954 sg13g2_dlygate4sd3_1
Xhold346 _0158_ VPWR VGND net965 sg13g2_dlygate4sd3_1
Xhold368 _0364_ VPWR VGND net987 sg13g2_dlygate4sd3_1
Xhold357 mydesign.pe_inputs\[13\] VPWR VGND net976 sg13g2_dlygate4sd3_1
X_4465_ _1389_ _1387_ _1388_ VPWR VGND sg13g2_xnor2_1
X_4396_ _1319_ VPWR _1323_ VGND _1305_ _1320_ sg13g2_o21ai_1
X_3416_ _0407_ VPWR _0461_ VGND net504 _0458_ sg13g2_o21ai_1
Xhold379 mydesign.accum\[110\] VPWR VGND net998 sg13g2_dlygate4sd3_1
X_3347_ net454 _2598_ net744 _0400_ VPWR VGND _2603_ sg13g2_nand4_1
X_6135_ net320 VGND VPWR _0361_ mydesign.weights\[0\]\[17\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_6066_ net194 VGND VPWR net696 mydesign.weights\[2\]\[8\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_3278_ _2682_ VPWR _0036_ VGND _2517_ _2678_ sg13g2_o21ai_1
X_5017_ _1869_ VPWR _1870_ VGND net591 net1019 sg13g2_o21ai_1
XFILLER_26_401 VPWR VGND sg13g2_decap_8
XFILLER_42_905 VPWR VGND sg13g2_decap_8
XFILLER_14_629 VPWR VGND sg13g2_fill_2
XFILLER_41_448 VPWR VGND sg13g2_fill_2
XFILLER_13_117 VPWR VGND sg13g2_decap_4
XFILLER_13_128 VPWR VGND sg13g2_fill_2
X_5919_ net319 VGND VPWR _0145_ mydesign.accum\[101\] clknet_leaf_45_clk sg13g2_dfrbpq_2
XFILLER_10_879 VPWR VGND sg13g2_decap_8
XFILLER_1_522 VPWR VGND sg13g2_fill_2
XFILLER_27_1011 VPWR VGND sg13g2_decap_8
XFILLER_18_946 VPWR VGND sg13g2_decap_8
XFILLER_45_765 VPWR VGND sg13g2_decap_8
XFILLER_33_938 VPWR VGND sg13g2_decap_8
XFILLER_41_993 VPWR VGND sg13g2_decap_8
XFILLER_40_470 VPWR VGND sg13g2_decap_8
XFILLER_8_110 VPWR VGND sg13g2_fill_1
XFILLER_34_1026 VPWR VGND sg13g2_fill_2
XFILLER_8_187 VPWR VGND sg13g2_fill_1
XFILLER_5_883 VPWR VGND sg13g2_decap_4
X_4250_ _1194_ mydesign.pe_weights\[56\] mydesign.pe_inputs\[46\] VPWR VGND sg13g2_nand2_1
X_4181_ VGND VPWR net569 _1137_ _0160_ _1138_ sg13g2_a21oi_1
X_3201_ _2633_ _2632_ VPWR VGND _2605_ sg13g2_nand2b_2
X_3132_ VPWR _2573_ net999 VGND sg13g2_inv_1
XFILLER_35_220 VPWR VGND sg13g2_fill_2
X_3965_ _0914_ mydesign.pe_inputs\[53\] _0942_ VPWR VGND sg13g2_nor2b_1
X_5704_ _2479_ VPWR _0342_ VGND net599 _2476_ sg13g2_o21ai_1
X_3896_ _0884_ VPWR _0885_ VGND _0864_ _0866_ sg13g2_o21ai_1
XFILLER_31_470 VPWR VGND sg13g2_decap_8
XFILLER_32_971 VPWR VGND sg13g2_decap_8
X_5635_ _2425_ _2404_ _2424_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_809 VPWR VGND sg13g2_decap_8
X_5566_ _2360_ VPWR _0323_ VGND net597 _2355_ sg13g2_o21ai_1
Xhold110 mydesign.accum\[8\] VPWR VGND net729 sg13g2_dlygate4sd3_1
Xhold121 _0172_ VPWR VGND net740 sg13g2_dlygate4sd3_1
X_4517_ _1427_ _1424_ _1429_ VPWR VGND sg13g2_xor2_1
Xhold132 mydesign.weights\[0\]\[19\] VPWR VGND net751 sg13g2_dlygate4sd3_1
X_5497_ mydesign.pe_inputs\[10\] net525 mydesign.accum\[12\] _2299_ VPWR VGND sg13g2_nand3_1
Xhold143 mydesign.inputs\[1\]\[12\] VPWR VGND net762 sg13g2_dlygate4sd3_1
Xhold176 mydesign.inputs\[1\]\[20\] VPWR VGND net795 sg13g2_dlygate4sd3_1
Xhold165 mydesign.weights\[0\]\[14\] VPWR VGND net784 sg13g2_dlygate4sd3_1
X_4448_ _1351_ VPWR _1373_ VGND _1344_ _1352_ sg13g2_o21ai_1
Xhold154 mydesign.accum\[27\] VPWR VGND net773 sg13g2_dlygate4sd3_1
Xhold187 mydesign.accum\[94\] VPWR VGND net806 sg13g2_dlygate4sd3_1
Xhold198 _0271_ VPWR VGND net817 sg13g2_dlygate4sd3_1
Xfanout612 net613 net612 VPWR VGND sg13g2_buf_8
Xfanout623 net627 net623 VPWR VGND sg13g2_buf_8
Xfanout601 _2627_ net601 VPWR VGND sg13g2_buf_8
X_4379_ VGND VPWR net573 _1306_ _0189_ _1307_ sg13g2_a21oi_1
Xfanout634 net636 net634 VPWR VGND sg13g2_buf_8
X_6118_ net92 VGND VPWR _0344_ mydesign.weights\[1\]\[8\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_6049_ net262 VGND VPWR _0275_ mydesign.accum\[35\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_2_1013 VPWR VGND sg13g2_decap_8
XFILLER_37_57 VPWR VGND sg13g2_decap_8
XFILLER_27_776 VPWR VGND sg13g2_decap_8
XFILLER_10_632 VPWR VGND sg13g2_decap_8
XFILLER_6_669 VPWR VGND sg13g2_decap_4
XFILLER_5_124 VPWR VGND sg13g2_decap_4
XFILLER_1_363 VPWR VGND sg13g2_fill_2
XFILLER_49_334 VPWR VGND sg13g2_fill_1
XFILLER_37_518 VPWR VGND sg13g2_decap_4
XFILLER_17_220 VPWR VGND sg13g2_fill_1
X_6130__364 VPWR VGND net364 sg13g2_tiehi
XFILLER_17_253 VPWR VGND sg13g2_fill_2
XFILLER_32_223 VPWR VGND sg13g2_fill_2
XFILLER_33_724 VPWR VGND sg13g2_fill_1
X_3750_ _0757_ VPWR _0758_ VGND _0725_ _0726_ sg13g2_o21ai_1
XFILLER_32_278 VPWR VGND sg13g2_fill_1
X_3681_ _0692_ mydesign.accum\[115\] net540 _0658_ VPWR VGND sg13g2_and3_1
X_5420_ _2232_ _2218_ _2215_ VPWR VGND sg13g2_nand2b_1
X_5351_ VGND VPWR net591 _2165_ _0302_ _2166_ sg13g2_a21oi_1
X_4302_ _1244_ _1242_ _1243_ VPWR VGND sg13g2_nand2_1
X_5282_ VGND VPWR net565 _2109_ _0289_ _2110_ sg13g2_a21oi_1
X_4233_ VGND VPWR _2565_ net448 _0170_ _1180_ sg13g2_a21oi_1
X_4164_ _1122_ _1104_ _1102_ VPWR VGND sg13g2_nand2b_1
X_4095_ net626 VPWR _1062_ VGND net489 _1061_ sg13g2_o21ai_1
X_3115_ VPWR _2556_ net538 VGND sg13g2_inv_1
X_4997_ _1849_ VPWR _1851_ VGND _1828_ _1830_ sg13g2_o21ai_1
X_3948_ VGND VPWR _2554_ net486 _0138_ _0927_ sg13g2_a21oi_1
XFILLER_32_790 VPWR VGND sg13g2_decap_8
X_3879_ _0869_ _0856_ _0867_ VPWR VGND sg13g2_xnor2_1
X_5618_ _2408_ mydesign.pe_inputs\[5\] mydesign.pe_weights\[19\] VPWR VGND sg13g2_nand2_1
XFILLER_20_996 VPWR VGND sg13g2_decap_8
XFILLER_3_606 VPWR VGND sg13g2_decap_4
X_5903__347 VPWR VGND net347 sg13g2_tiehi
X_5549_ _2348_ _2342_ _2345_ VPWR VGND sg13g2_nand2_1
XFILLER_3_639 VPWR VGND sg13g2_fill_2
X_6123__48 VPWR VGND net48 sg13g2_tiehi
Xfanout431 _2697_ net431 VPWR VGND sg13g2_buf_8
Xfanout475 net477 net475 VPWR VGND sg13g2_buf_8
Xfanout442 net446 net442 VPWR VGND sg13g2_buf_8
Xfanout464 net466 net464 VPWR VGND sg13g2_buf_8
Xfanout453 _2601_ net453 VPWR VGND sg13g2_buf_8
XFILLER_47_838 VPWR VGND sg13g2_decap_8
XFILLER_48_89 VPWR VGND sg13g2_fill_1
Xfanout497 _2587_ net497 VPWR VGND sg13g2_buf_8
XFILLER_19_507 VPWR VGND sg13g2_fill_2
Xfanout486 net490 net486 VPWR VGND sg13g2_buf_8
XFILLER_42_532 VPWR VGND sg13g2_decap_8
X_5947__263 VPWR VGND net263 sg13g2_tiehi
XFILLER_7_967 VPWR VGND sg13g2_decap_8
XFILLER_11_996 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_fill_1
XFILLER_9_1019 VPWR VGND sg13g2_decap_8
XFILLER_38_827 VPWR VGND sg13g2_decap_8
XFILLER_37_315 VPWR VGND sg13g2_fill_2
X_4920_ VGND VPWR _2536_ net445 _0256_ _1781_ sg13g2_a21oi_1
XFILLER_18_584 VPWR VGND sg13g2_decap_4
XFILLER_18_595 VPWR VGND sg13g2_decap_4
XFILLER_33_510 VPWR VGND sg13g2_decap_4
X_4851_ mydesign.pe_inputs\[30\] net533 mydesign.accum\[53\] _1728_ VPWR VGND sg13g2_a21o_1
X_3802_ VGND VPWR _2557_ net491 _0122_ _0797_ sg13g2_a21oi_1
X_4782_ _1661_ _1662_ _1663_ VPWR VGND sg13g2_nor2b_1
X_3733_ _0742_ _0721_ _0741_ VPWR VGND sg13g2_nand2_1
X_3664_ _0674_ _0675_ _0676_ VPWR VGND sg13g2_nor2_1
X_5403_ _2214_ _2213_ _2216_ VPWR VGND sg13g2_xor2_1
X_3595_ _0619_ _0616_ _0618_ VPWR VGND sg13g2_nand2_1
X_6137__304 VPWR VGND net304 sg13g2_tiehi
X_5334_ net481 VPWR _2151_ VGND net591 net1029 sg13g2_o21ai_1
X_5265_ VGND VPWR _2075_ _2091_ _2094_ _2090_ sg13g2_a21oi_1
X_4216_ _1171_ _1161_ _1170_ VPWR VGND sg13g2_xnor2_1
X_5196_ _2027_ _2028_ _2029_ VPWR VGND sg13g2_nor2_1
X_4147_ _1106_ _1081_ _1104_ _1105_ VPWR VGND sg13g2_and3_1
X_4078_ VGND VPWR _2571_ net488 _0148_ _1047_ sg13g2_a21oi_1
Xclkload2 clknet_3_3__leaf_clk clkload2/X VPWR VGND sg13g2_buf_8
XFILLER_20_771 VPWR VGND sg13g2_fill_1
XFILLER_4_948 VPWR VGND sg13g2_decap_8
XFILLER_3_469 VPWR VGND sg13g2_decap_4
XFILLER_47_635 VPWR VGND sg13g2_decap_8
XFILLER_43_830 VPWR VGND sg13g2_decap_8
XFILLER_15_521 VPWR VGND sg13g2_fill_2
XFILLER_28_893 VPWR VGND sg13g2_decap_8
XFILLER_15_543 VPWR VGND sg13g2_fill_1
X_6088__380 VPWR VGND net380 sg13g2_tiehi
XFILLER_30_568 VPWR VGND sg13g2_fill_2
X_3380_ VGND VPWR _0419_ _0427_ _0069_ _0428_ sg13g2_a21oi_1
XFILLER_3_992 VPWR VGND sg13g2_decap_8
X_5050_ VGND VPWR net734 _1894_ _0272_ _1895_ sg13g2_a21oi_1
X_4001_ _0967_ VPWR _0976_ VGND _0973_ _0974_ sg13g2_o21ai_1
XFILLER_38_635 VPWR VGND sg13g2_decap_8
X_5952_ net253 VGND VPWR _0178_ mydesign.accum\[86\] clknet_leaf_25_clk sg13g2_dfrbpq_2
XFILLER_19_882 VPWR VGND sg13g2_fill_1
XFILLER_25_318 VPWR VGND sg13g2_fill_2
X_4903_ net612 VPWR _1772_ VGND net858 _1767_ sg13g2_o21ai_1
XFILLER_34_863 VPWR VGND sg13g2_decap_4
X_5883_ net383 VGND VPWR _0109_ mydesign.accum\[117\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4834_ _1712_ _1705_ _1711_ VPWR VGND sg13g2_nand2_1
X_4765_ VGND VPWR _2545_ net447 _0231_ _1651_ sg13g2_a21oi_1
X_3716_ VGND VPWR _0687_ _0706_ _0726_ _0705_ sg13g2_a21oi_1
X_4696_ _1591_ _1571_ _1590_ VPWR VGND sg13g2_xnor2_1
X_5822__120 VPWR VGND net120 sg13g2_tiehi
XFILLER_20_49 VPWR VGND sg13g2_fill_1
X_3647_ _0661_ net577 _0660_ VPWR VGND sg13g2_nand2_1
X_3578_ _0600_ _0602_ _0603_ VPWR VGND sg13g2_nor2_1
XFILLER_1_929 VPWR VGND sg13g2_decap_8
X_5317_ VGND VPWR _2523_ net493 _0297_ _2137_ sg13g2_a21oi_1
Xhold14 mydesign.inputs\[2\]\[9\] VPWR VGND net420 sg13g2_dlygate4sd3_1
Xhold25 mydesign.inputs\[3\]\[13\] VPWR VGND net644 sg13g2_dlygate4sd3_1
Xhold47 mydesign.inputs\[3\]\[15\] VPWR VGND net666 sg13g2_dlygate4sd3_1
X_5248_ _2078_ mydesign.pe_weights\[29\] _2020_ VPWR VGND sg13g2_nand2_1
Xhold36 mydesign.inputs\[2\]\[4\] VPWR VGND net655 sg13g2_dlygate4sd3_1
X_5179_ _2014_ VPWR _2015_ VGND _2012_ _2013_ sg13g2_o21ai_1
Xhold69 mydesign.accum\[104\] VPWR VGND net688 sg13g2_dlygate4sd3_1
Xhold58 mydesign.weights\[2\]\[16\] VPWR VGND net677 sg13g2_dlygate4sd3_1
XFILLER_44_638 VPWR VGND sg13g2_decap_8
XFILLER_24_362 VPWR VGND sg13g2_fill_1
XFILLER_12_535 VPWR VGND sg13g2_fill_1
XFILLER_4_701 VPWR VGND sg13g2_fill_1
XFILLER_48_944 VPWR VGND sg13g2_decap_8
X_6051__254 VPWR VGND net254 sg13g2_tiehi
XFILLER_47_498 VPWR VGND sg13g2_fill_1
XFILLER_35_627 VPWR VGND sg13g2_decap_8
XFILLER_34_126 VPWR VGND sg13g2_fill_1
XFILLER_16_896 VPWR VGND sg13g2_fill_2
X_4550_ _1443_ VPWR _1460_ VGND _1442_ _1445_ sg13g2_o21ai_1
XFILLER_7_561 VPWR VGND sg13g2_fill_1
X_4481_ _1403_ net646 _1402_ VPWR VGND sg13g2_nand2_1
X_3501_ net455 _0520_ mydesign.accum\[121\] _0530_ VPWR VGND sg13g2_nand3_1
X_3432_ _0405_ VPWR _0476_ VGND net509 _0473_ sg13g2_o21ai_1
X_3363_ _0412_ VPWR _0413_ VGND net507 _0409_ sg13g2_o21ai_1
X_5102_ _1944_ mydesign.pe_weights\[35\] mydesign.pe_inputs\[21\] VPWR VGND sg13g2_nand2_1
XFILLER_39_900 VPWR VGND sg13g2_decap_8
X_6082_ net52 VGND VPWR net1066 mydesign.pe_inputs\[4\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3294_ VGND VPWR net608 _2690_ _2689_ net605 sg13g2_a21oi_2
Xheichips25_template_16 VPWR VGND uio_out[1] sg13g2_tielo
X_5033_ _1881_ VPWR _1884_ VGND _1862_ _1878_ sg13g2_o21ai_1
XFILLER_39_977 VPWR VGND sg13g2_decap_8
X_5935_ net287 VGND VPWR _0161_ mydesign.accum\[93\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_5866_ net41 VGND VPWR _0092_ mydesign.accum\[124\] clknet_leaf_16_clk sg13g2_dfrbpq_2
XFILLER_40_129 VPWR VGND sg13g2_fill_1
XFILLER_33_170 VPWR VGND sg13g2_fill_1
X_4817_ _1696_ _1673_ _1695_ VPWR VGND sg13g2_nand2_1
X_5797_ net153 VGND VPWR _0023_ mydesign.inputs\[1\]\[10\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_22_899 VPWR VGND sg13g2_fill_1
X_4748_ _1640_ _1630_ _1639_ VPWR VGND sg13g2_xnor2_1
X_4679_ _1574_ mydesign.pe_weights\[45\] _1531_ VPWR VGND sg13g2_nand2b_1
Xoutput15 net15 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_737 VPWR VGND sg13g2_fill_1
XFILLER_5_1000 VPWR VGND sg13g2_decap_8
XFILLER_29_454 VPWR VGND sg13g2_fill_2
XFILLER_45_947 VPWR VGND sg13g2_decap_8
XFILLER_16_126 VPWR VGND sg13g2_fill_1
XFILLER_16_148 VPWR VGND sg13g2_fill_2
XFILLER_31_107 VPWR VGND sg13g2_fill_1
XFILLER_13_844 VPWR VGND sg13g2_fill_1
X_6010__50 VPWR VGND net50 sg13g2_tiehi
XFILLER_21_92 VPWR VGND sg13g2_decap_4
XFILLER_39_207 VPWR VGND sg13g2_decap_8
XFILLER_48_741 VPWR VGND sg13g2_decap_8
XFILLER_35_402 VPWR VGND sg13g2_decap_8
XFILLER_36_958 VPWR VGND sg13g2_decap_8
X_5812__130 VPWR VGND net130 sg13g2_tiehi
X_3981_ _0949_ _0956_ _0957_ VPWR VGND sg13g2_nor2b_1
X_5720_ net771 _2485_ _2489_ _0348_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_42_clk clknet_3_4__leaf_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
X_5651_ _2438_ _2428_ _2440_ VPWR VGND sg13g2_xor2_1
XFILLER_31_674 VPWR VGND sg13g2_decap_8
XFILLER_31_685 VPWR VGND sg13g2_fill_1
X_4602_ _1506_ VPWR _1509_ VGND _1489_ _1502_ sg13g2_o21ai_1
X_5582_ _2365_ VPWR _2374_ VGND _2363_ _2366_ sg13g2_o21ai_1
XFILLER_30_195 VPWR VGND sg13g2_decap_8
XFILLER_8_892 VPWR VGND sg13g2_fill_1
XFILLER_8_881 VPWR VGND sg13g2_fill_1
X_4533_ net532 net537 mydesign.accum\[67\] _1444_ VPWR VGND sg13g2_a21o_1
Xhold314 mydesign.accum\[84\] VPWR VGND net933 sg13g2_dlygate4sd3_1
Xhold325 mydesign.accum\[102\] VPWR VGND net944 sg13g2_dlygate4sd3_1
Xhold303 _0262_ VPWR VGND net922 sg13g2_dlygate4sd3_1
Xhold369 mydesign.pe_weights\[58\] VPWR VGND net988 sg13g2_dlygate4sd3_1
Xhold347 mydesign.pe_inputs\[37\] VPWR VGND net966 sg13g2_dlygate4sd3_1
Xhold336 _0285_ VPWR VGND net955 sg13g2_dlygate4sd3_1
X_4464_ _1388_ _1374_ _1371_ VPWR VGND sg13g2_nand2b_1
Xhold358 mydesign.accum\[79\] VPWR VGND net977 sg13g2_dlygate4sd3_1
X_4395_ VGND VPWR net575 _1321_ _0190_ _1322_ sg13g2_a21oi_1
X_3415_ VGND VPWR net890 net512 _0460_ _0459_ sg13g2_a21oi_1
X_3346_ VGND VPWR net454 _2603_ _0399_ net744 sg13g2_a21oi_1
X_6134_ net328 VGND VPWR _0360_ mydesign.weights\[0\]\[16\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_6065_ net198 VGND VPWR _0291_ mydesign.accum\[31\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_3277_ net616 _2678_ net736 _2682_ VPWR VGND sg13g2_nand3_1
X_5016_ net591 VPWR _1869_ VGND _1867_ _1868_ sg13g2_o21ai_1
XFILLER_38_240 VPWR VGND sg13g2_fill_2
XFILLER_27_969 VPWR VGND sg13g2_decap_8
XFILLER_26_479 VPWR VGND sg13g2_fill_1
XFILLER_41_416 VPWR VGND sg13g2_decap_8
X_5918_ net321 VGND VPWR _0144_ mydesign.accum\[100\] clknet_leaf_46_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_33_clk clknet_3_7__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
XFILLER_22_652 VPWR VGND sg13g2_fill_2
X_6106__228 VPWR VGND net228 sg13g2_tiehi
XFILLER_21_140 VPWR VGND sg13g2_fill_2
X_5849_ net71 VGND VPWR net1085 net15 clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_10_847 VPWR VGND sg13g2_decap_8
XFILLER_1_534 VPWR VGND sg13g2_fill_1
XFILLER_17_402 VPWR VGND sg13g2_decap_8
XFILLER_29_262 VPWR VGND sg13g2_fill_1
XFILLER_45_744 VPWR VGND sg13g2_decap_8
XFILLER_17_424 VPWR VGND sg13g2_fill_2
XFILLER_29_284 VPWR VGND sg13g2_fill_2
XFILLER_33_917 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_24_clk clknet_3_6__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_34_1005 VPWR VGND sg13g2_decap_8
XFILLER_41_972 VPWR VGND sg13g2_decap_8
XFILLER_12_151 VPWR VGND sg13g2_decap_8
XFILLER_8_144 VPWR VGND sg13g2_fill_2
XFILLER_4_394 VPWR VGND sg13g2_fill_2
X_4180_ net468 VPWR _1138_ VGND net569 net997 sg13g2_o21ai_1
X_5957__243 VPWR VGND net243 sg13g2_tiehi
X_3200_ _2606_ _2622_ _2632_ VPWR VGND sg13g2_nor2_2
X_3131_ VPWR _2572_ mydesign.accum\[94\] VGND sg13g2_inv_1
Xclkbuf_leaf_15_clk clknet_3_2__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_3964_ VGND VPWR _0941_ _0940_ _0939_ sg13g2_or2_1
XFILLER_32_950 VPWR VGND sg13g2_decap_8
X_5703_ net705 _2476_ net613 _2479_ VPWR VGND sg13g2_nand3_1
X_3895_ _0882_ _0881_ _0884_ VPWR VGND sg13g2_xor2_1
X_5634_ _2424_ _2407_ _2422_ VPWR VGND sg13g2_xnor2_1
Xhold100 mydesign.inputs\[3\]\[3\] VPWR VGND net719 sg13g2_dlygate4sd3_1
X_5565_ _2360_ net680 _2356_ VPWR VGND sg13g2_nand2_1
X_4516_ _1424_ _1427_ _1428_ VPWR VGND sg13g2_nor2_1
Xhold122 mydesign.weights\[2\]\[6\] VPWR VGND net741 sg13g2_dlygate4sd3_1
Xhold133 mydesign.weights\[2\]\[7\] VPWR VGND net752 sg13g2_dlygate4sd3_1
Xhold111 _0312_ VPWR VGND net730 sg13g2_dlygate4sd3_1
X_5496_ _2298_ mydesign.pe_inputs\[9\] mydesign.pe_weights\[23\] VPWR VGND sg13g2_nand2_1
Xhold144 mydesign.weights\[1\]\[15\] VPWR VGND net763 sg13g2_dlygate4sd3_1
Xhold166 mydesign.inputs\[0\]\[22\] VPWR VGND net785 sg13g2_dlygate4sd3_1
X_4447_ _1370_ _1369_ _1372_ VPWR VGND sg13g2_xor2_1
Xhold155 mydesign.weights\[1\]\[9\] VPWR VGND net774 sg13g2_dlygate4sd3_1
Xhold177 mydesign.inputs\[1\]\[16\] VPWR VGND net796 sg13g2_dlygate4sd3_1
Xfanout613 net619 net613 VPWR VGND sg13g2_buf_8
Xhold188 mydesign.weights\[2\]\[13\] VPWR VGND net807 sg13g2_dlygate4sd3_1
Xfanout602 _2627_ net602 VPWR VGND sg13g2_buf_8
Xfanout624 net627 net624 VPWR VGND sg13g2_buf_8
Xhold199 mydesign.accum\[57\] VPWR VGND net818 sg13g2_dlygate4sd3_1
X_6117_ net100 VGND VPWR net732 mydesign.weights\[3\]\[3\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_4378_ net478 VPWR _1307_ VGND net573 net875 sg13g2_o21ai_1
Xfanout635 net636 net635 VPWR VGND sg13g2_buf_2
X_3329_ VGND VPWR net563 _2600_ _0386_ _0385_ sg13g2_a21oi_1
XFILLER_37_14 VPWR VGND sg13g2_fill_1
X_6048_ net266 VGND VPWR net914 mydesign.accum\[34\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_23_994 VPWR VGND sg13g2_decap_8
XFILLER_10_688 VPWR VGND sg13g2_fill_2
X_6126__24 VPWR VGND net24 sg13g2_tiehi
XFILLER_5_169 VPWR VGND sg13g2_fill_2
XFILLER_5_158 VPWR VGND sg13g2_decap_8
XFILLER_1_320 VPWR VGND sg13g2_fill_2
XFILLER_18_788 VPWR VGND sg13g2_fill_2
XFILLER_17_265 VPWR VGND sg13g2_fill_2
XFILLER_32_202 VPWR VGND sg13g2_decap_8
XFILLER_33_714 VPWR VGND sg13g2_decap_4
X_3680_ _0691_ mydesign.pe_inputs\[61\] _0653_ VPWR VGND sg13g2_nand2_1
X_5350_ net481 VPWR _2166_ VGND net590 net1020 sg13g2_o21ai_1
X_4301_ _1222_ VPWR _1243_ VGND _1211_ _1223_ sg13g2_o21ai_1
X_5281_ net465 VPWR _2110_ VGND net565 net890 sg13g2_o21ai_1
X_4232_ net631 VPWR _1180_ VGND net813 net448 sg13g2_o21ai_1
Xclkbuf_leaf_4_clk clknet_3_0__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_4163_ _1121_ mydesign.pe_weights\[61\] _1061_ VPWR VGND sg13g2_nand2_1
X_4094_ _0639_ net800 _1060_ _1061_ VPWR VGND sg13g2_a21o_2
X_3114_ _2555_ net872 VPWR VGND sg13g2_inv_2
X_4996_ _1828_ _1830_ _1849_ _1850_ VPWR VGND sg13g2_or3_1
XFILLER_24_769 VPWR VGND sg13g2_decap_8
X_3947_ net628 VPWR _0927_ VGND net486 _0926_ sg13g2_o21ai_1
XFILLER_11_419 VPWR VGND sg13g2_decap_4
X_3878_ _0868_ _0856_ _0867_ VPWR VGND sg13g2_nand2_1
XFILLER_20_975 VPWR VGND sg13g2_decap_8
X_5617_ _2401_ VPWR _2407_ VGND _2387_ _2402_ sg13g2_o21ai_1
X_5548_ VGND VPWR net592 _2346_ _0318_ _2347_ sg13g2_a21oi_1
X_5479_ _2282_ _2280_ _2281_ VPWR VGND sg13g2_nand2_1
Xfanout432 _2608_ net432 VPWR VGND sg13g2_buf_8
Xfanout454 _2596_ net454 VPWR VGND sg13g2_buf_8
Xfanout443 net446 net443 VPWR VGND sg13g2_buf_1
Xfanout465 net466 net465 VPWR VGND sg13g2_buf_8
XFILLER_47_817 VPWR VGND sg13g2_decap_8
Xfanout498 _2587_ net498 VPWR VGND sg13g2_buf_8
Xfanout476 net477 net476 VPWR VGND sg13g2_buf_2
Xfanout487 net490 net487 VPWR VGND sg13g2_buf_8
XFILLER_27_530 VPWR VGND sg13g2_fill_1
XFILLER_15_769 VPWR VGND sg13g2_decap_4
X_6047__270 VPWR VGND net270 sg13g2_tiehi
XFILLER_11_975 VPWR VGND sg13g2_decap_8
XFILLER_49_154 VPWR VGND sg13g2_decap_4
XFILLER_38_817 VPWR VGND sg13g2_decap_4
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_46_894 VPWR VGND sg13g2_decap_8
X_4850_ net533 mydesign.pe_inputs\[30\] mydesign.accum\[53\] _1727_ VPWR VGND sg13g2_nand3_1
X_3801_ net628 VPWR _0797_ VGND net491 _0796_ sg13g2_o21ai_1
X_4781_ _1660_ VPWR _1662_ VGND _1658_ _1659_ sg13g2_o21ai_1
X_3732_ _0741_ _0731_ _0739_ VPWR VGND sg13g2_xnor2_1
X_5809__135 VPWR VGND net135 sg13g2_tiehi
X_6096__308 VPWR VGND net308 sg13g2_tiehi
X_3663_ VGND VPWR net540 _0653_ _0675_ mydesign.accum\[114\] sg13g2_a21oi_1
X_5402_ _2213_ _2214_ _2215_ VPWR VGND sg13g2_and2_1
X_3594_ _0526_ _0512_ mydesign.accum\[126\] _0618_ VPWR VGND sg13g2_a21o_1
X_5333_ _2148_ _2147_ _2150_ VPWR VGND sg13g2_xor2_1
X_5264_ VGND VPWR net565 _2092_ _0288_ _2093_ sg13g2_a21oi_1
X_4215_ _1169_ net948 _1170_ VPWR VGND sg13g2_xor2_1
X_5195_ _2028_ net891 _2010_ VPWR VGND sg13g2_nand2_1
X_4146_ _1101_ VPWR _1105_ VGND _1102_ _1103_ sg13g2_o21ai_1
X_4077_ net626 VPWR _1047_ VGND net489 _1046_ sg13g2_o21ai_1
XFILLER_43_308 VPWR VGND sg13g2_fill_2
X_4979_ _1833_ mydesign.pe_weights\[37\] mydesign.pe_inputs\[27\] VPWR VGND sg13g2_nand2_1
Xclkload3 clknet_3_5__leaf_clk clkload3/X VPWR VGND sg13g2_buf_8
XFILLER_47_614 VPWR VGND sg13g2_decap_8
XFILLER_46_146 VPWR VGND sg13g2_decap_8
XFILLER_27_371 VPWR VGND sg13g2_decap_8
XFILLER_43_886 VPWR VGND sg13g2_decap_8
XFILLER_24_70 VPWR VGND sg13g2_fill_1
XFILLER_24_92 VPWR VGND sg13g2_decap_4
XFILLER_7_798 VPWR VGND sg13g2_fill_2
XFILLER_6_286 VPWR VGND sg13g2_fill_2
XFILLER_3_971 VPWR VGND sg13g2_decap_8
XFILLER_2_470 VPWR VGND sg13g2_decap_8
X_4000_ _0967_ _0973_ _0974_ _0975_ VPWR VGND sg13g2_or3_1
XFILLER_38_658 VPWR VGND sg13g2_fill_2
XFILLER_37_157 VPWR VGND sg13g2_fill_1
X_5951_ net255 VGND VPWR _0177_ mydesign.accum\[85\] clknet_leaf_25_clk sg13g2_dfrbpq_2
XFILLER_46_691 VPWR VGND sg13g2_decap_8
X_4902_ _1771_ net2 _1768_ VPWR VGND sg13g2_nand2_2
XFILLER_34_886 VPWR VGND sg13g2_decap_8
X_5882_ net385 VGND VPWR _0108_ mydesign.accum\[116\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_4833_ _1709_ _1706_ _1711_ VPWR VGND sg13g2_xor2_1
X_4764_ net637 VPWR _1651_ VGND mydesign.pe_inputs\[27\] net447 sg13g2_o21ai_1
X_3715_ _0725_ _0724_ VPWR VGND _0723_ sg13g2_nand2b_2
X_4695_ _1590_ _1572_ _1588_ VPWR VGND sg13g2_xnor2_1
X_3646_ net540 _0643_ _0660_ VPWR VGND sg13g2_and2_1
X_3577_ _0602_ mydesign.accum\[125\] _0601_ VPWR VGND sg13g2_xnor2_1
XFILLER_1_908 VPWR VGND sg13g2_decap_8
XFILLER_0_407 VPWR VGND sg13g2_decap_8
X_5316_ net634 VPWR _2137_ VGND net976 net493 sg13g2_o21ai_1
X_5247_ _2077_ _2061_ _2063_ VPWR VGND sg13g2_nand2_1
Xhold37 mydesign.weights\[2\]\[11\] VPWR VGND net656 sg13g2_dlygate4sd3_1
Xhold15 _0014_ VPWR VGND net421 sg13g2_dlygate4sd3_1
Xhold26 mydesign.weights\[1\]\[18\] VPWR VGND net645 sg13g2_dlygate4sd3_1
X_5178_ _2014_ _0395_ mydesign.inputs\[3\]\[14\] net454 mydesign.inputs\[3\]\[2\]
+ VPWR VGND sg13g2_a22oi_1
Xhold59 _0009_ VPWR VGND net678 sg13g2_dlygate4sd3_1
Xhold48 mydesign.inputs\[2\]\[10\] VPWR VGND net667 sg13g2_dlygate4sd3_1
X_4129_ _1089_ _1088_ _1080_ VPWR VGND sg13g2_nand2b_1
XFILLER_45_69 VPWR VGND sg13g2_fill_1
XFILLER_40_834 VPWR VGND sg13g2_decap_4
XFILLER_40_889 VPWR VGND sg13g2_decap_8
XFILLER_20_580 VPWR VGND sg13g2_decap_4
XFILLER_4_746 VPWR VGND sg13g2_decap_8
XFILLER_3_278 VPWR VGND sg13g2_fill_2
X_5797__153 VPWR VGND net153 sg13g2_tiehi
XFILLER_48_923 VPWR VGND sg13g2_decap_8
X_5916__325 VPWR VGND net325 sg13g2_tiehi
XFILLER_0_985 VPWR VGND sg13g2_decap_8
XFILLER_19_113 VPWR VGND sg13g2_fill_2
XFILLER_34_105 VPWR VGND sg13g2_fill_2
XFILLER_43_650 VPWR VGND sg13g2_decap_8
XFILLER_15_341 VPWR VGND sg13g2_decap_4
XFILLER_43_694 VPWR VGND sg13g2_decap_8
XFILLER_15_385 VPWR VGND sg13g2_fill_2
XFILLER_30_311 VPWR VGND sg13g2_decap_4
XFILLER_31_834 VPWR VGND sg13g2_fill_2
XFILLER_30_344 VPWR VGND sg13g2_decap_4
XFILLER_30_388 VPWR VGND sg13g2_fill_2
XFILLER_7_551 VPWR VGND sg13g2_fill_2
X_3500_ VGND VPWR net721 _0528_ _0088_ _0529_ sg13g2_a21oi_1
X_4480_ net618 _1401_ _1402_ VPWR VGND sg13g2_and2_1
X_3431_ VGND VPWR mydesign.accum\[22\] net516 _0475_ _0474_ sg13g2_a21oi_1
X_3362_ net755 net834 _0412_ VPWR VGND sg13g2_nor2b_2
X_5101_ _1926_ VPWR _1943_ VGND _1925_ _1928_ sg13g2_o21ai_1
X_6081_ net60 VGND VPWR _0307_ mydesign.accum\[23\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_3293_ net596 _2688_ _2689_ VPWR VGND sg13g2_nor2_1
Xheichips25_template_17 VPWR VGND uio_out[2] sg13g2_tielo
X_5032_ _1882_ _1883_ _0266_ VPWR VGND sg13g2_nor2_1
XFILLER_39_956 VPWR VGND sg13g2_decap_8
XFILLER_38_477 VPWR VGND sg13g2_fill_1
XFILLER_25_127 VPWR VGND sg13g2_fill_1
X_5934_ net289 VGND VPWR _0160_ mydesign.accum\[92\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_5967__223 VPWR VGND net223 sg13g2_tiehi
X_5865_ net43 VGND VPWR _0091_ mydesign.accum\[123\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_4816_ _1693_ _1686_ _1695_ VPWR VGND sg13g2_xor2_1
X_5796_ net154 VGND VPWR _0022_ mydesign.inputs\[1\]\[9\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_4747_ _1637_ _1623_ _1639_ VPWR VGND sg13g2_xor2_1
X_4678_ _1573_ mydesign.pe_weights\[44\] _1537_ VPWR VGND sg13g2_nand2_1
X_3629_ _0646_ net461 mydesign.weights\[1\]\[21\] net495 mydesign.weights\[1\]\[17\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_0_259 VPWR VGND sg13g2_fill_2
XFILLER_0_248 VPWR VGND sg13g2_decap_8
XFILLER_29_444 VPWR VGND sg13g2_fill_2
XFILLER_45_926 VPWR VGND sg13g2_decap_8
XFILLER_40_675 VPWR VGND sg13g2_decap_4
XFILLER_4_510 VPWR VGND sg13g2_fill_1
X_5881__387 VPWR VGND net387 sg13g2_tiehi
XFILLER_4_532 VPWR VGND sg13g2_fill_1
X_6092__344 VPWR VGND net344 sg13g2_tiehi
XFILLER_48_720 VPWR VGND sg13g2_decap_8
XFILLER_0_760 VPWR VGND sg13g2_fill_2
XFILLER_0_782 VPWR VGND sg13g2_decap_8
XFILLER_48_797 VPWR VGND sg13g2_decap_8
XFILLER_36_937 VPWR VGND sg13g2_decap_8
X_3980_ _0956_ _0938_ _0955_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_609 VPWR VGND sg13g2_fill_1
XFILLER_44_981 VPWR VGND sg13g2_decap_8
XFILLER_16_694 VPWR VGND sg13g2_decap_8
X_5650_ _2439_ _2428_ _2438_ VPWR VGND sg13g2_nand2_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_30_130 VPWR VGND sg13g2_decap_8
X_4601_ _1507_ _1508_ _0210_ VPWR VGND sg13g2_nor2_1
X_5581_ _2373_ mydesign.pe_inputs\[4\] net1017 VPWR VGND sg13g2_nand2_1
X_4532_ net537 net532 mydesign.accum\[67\] _1443_ VPWR VGND sg13g2_nand3_1
XFILLER_11_1017 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
Xhold315 mydesign.pe_inputs\[9\] VPWR VGND net934 sg13g2_dlygate4sd3_1
X_4463_ _1387_ _1386_ _1385_ VPWR VGND sg13g2_nand2b_1
Xhold304 mydesign.accum\[26\] VPWR VGND net923 sg13g2_dlygate4sd3_1
Xhold326 mydesign.accum\[30\] VPWR VGND net945 sg13g2_dlygate4sd3_1
Xhold337 mydesign.pe_inputs\[47\] VPWR VGND net956 sg13g2_dlygate4sd3_1
Xhold359 mydesign.accum\[23\] VPWR VGND net978 sg13g2_dlygate4sd3_1
Xhold348 mydesign.accum\[99\] VPWR VGND net967 sg13g2_dlygate4sd3_1
X_3414_ net505 VPWR _0459_ VGND _2548_ net511 sg13g2_o21ai_1
X_4394_ net474 VPWR _1322_ VGND net575 net882 sg13g2_o21ai_1
X_3345_ VPWR VGND _0398_ net607 _0387_ _2586_ _0064_ _2604_ sg13g2_a221oi_1
X_6138__296 VPWR VGND net296 sg13g2_tiehi
X_6133_ net336 VGND VPWR _0359_ mydesign.weights\[0\]\[23\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3276_ _2681_ VPWR _0035_ VGND _2518_ _2678_ sg13g2_o21ai_1
X_6064_ net202 VGND VPWR _0290_ mydesign.accum\[30\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_5015_ VGND VPWR _1848_ _1851_ _1868_ _1866_ sg13g2_a21oi_1
XFILLER_27_948 VPWR VGND sg13g2_decap_8
X_5917_ net323 VGND VPWR _0143_ mydesign.accum\[99\] clknet_leaf_46_clk sg13g2_dfrbpq_2
XFILLER_35_992 VPWR VGND sg13g2_decap_8
XFILLER_22_686 VPWR VGND sg13g2_fill_1
X_5848_ net73 VGND VPWR _0074_ net14 clknet_leaf_7_clk sg13g2_dfrbpq_2
X_5787__163 VPWR VGND net163 sg13g2_tiehi
X_5779_ net175 VGND VPWR _0005_ mydesign.inputs\[0\]\[24\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_49_506 VPWR VGND sg13g2_decap_4
XFILLER_49_528 VPWR VGND sg13g2_decap_8
X_5794__156 VPWR VGND net156 sg13g2_tiehi
XFILLER_45_723 VPWR VGND sg13g2_decap_8
XFILLER_44_222 VPWR VGND sg13g2_fill_2
XFILLER_17_436 VPWR VGND sg13g2_fill_2
XFILLER_17_447 VPWR VGND sg13g2_fill_1
XFILLER_17_458 VPWR VGND sg13g2_fill_2
XFILLER_26_981 VPWR VGND sg13g2_decap_8
XFILLER_32_417 VPWR VGND sg13g2_decap_4
XFILLER_41_951 VPWR VGND sg13g2_decap_8
XFILLER_8_101 VPWR VGND sg13g2_fill_1
XFILLER_12_141 VPWR VGND sg13g2_decap_4
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_863 VPWR VGND sg13g2_fill_1
XFILLER_5_852 VPWR VGND sg13g2_fill_2
X_3130_ _2571_ net536 VPWR VGND sg13g2_inv_2
XFILLER_48_594 VPWR VGND sg13g2_decap_8
XFILLER_35_222 VPWR VGND sg13g2_fill_1
XFILLER_36_734 VPWR VGND sg13g2_decap_4
XFILLER_36_767 VPWR VGND sg13g2_decap_8
XFILLER_17_992 VPWR VGND sg13g2_decap_8
X_3963_ VGND VPWR mydesign.pe_inputs\[52\] _0919_ _0940_ mydesign.accum\[97\] sg13g2_a21oi_1
X_5702_ _2478_ VPWR _0341_ VGND net601 _2476_ sg13g2_o21ai_1
X_3894_ _0883_ _0881_ _0882_ VPWR VGND sg13g2_nand2_1
X_5633_ _2423_ _2407_ _2422_ VPWR VGND sg13g2_nand2_1
X_5564_ _2359_ VPWR _0322_ VGND net599 _2355_ sg13g2_o21ai_1
X_4515_ _1427_ _1425_ _1426_ VPWR VGND sg13g2_nand2_1
Xhold101 _0056_ VPWR VGND net720 sg13g2_dlygate4sd3_1
Xhold123 mydesign.inputs\[3\]\[1\] VPWR VGND net742 sg13g2_dlygate4sd3_1
Xhold112 mydesign.weights\[3\]\[3\] VPWR VGND net731 sg13g2_dlygate4sd3_1
Xhold134 _0004_ VPWR VGND net753 sg13g2_dlygate4sd3_1
X_5495_ _2280_ VPWR _2297_ VGND _2279_ _2282_ sg13g2_o21ai_1
Xhold156 mydesign.inputs\[1\]\[15\] VPWR VGND net775 sg13g2_dlygate4sd3_1
Xhold167 mydesign.inputs\[0\]\[13\] VPWR VGND net786 sg13g2_dlygate4sd3_1
X_4446_ _1369_ _1370_ _1371_ VPWR VGND sg13g2_and2_1
Xhold145 mydesign.weights\[1\]\[13\] VPWR VGND net764 sg13g2_dlygate4sd3_1
Xhold178 mydesign.inputs\[1\]\[14\] VPWR VGND net797 sg13g2_dlygate4sd3_1
Xhold189 mydesign.pe_weights\[60\] VPWR VGND net808 sg13g2_dlygate4sd3_1
X_4377_ _1304_ _1303_ _1306_ VPWR VGND sg13g2_xor2_1
Xfanout614 net615 net614 VPWR VGND sg13g2_buf_8
Xfanout603 _2625_ net603 VPWR VGND sg13g2_buf_8
X_6116_ net108 VGND VPWR net706 mydesign.weights\[3\]\[2\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_3328_ _0385_ _2692_ _0384_ VPWR VGND sg13g2_nand2_1
Xfanout636 net639 net636 VPWR VGND sg13g2_buf_8
Xfanout625 net626 net625 VPWR VGND sg13g2_buf_8
X_3259_ net797 _2669_ _2672_ _0027_ VPWR VGND sg13g2_mux2_1
X_6047_ net270 VGND VPWR net920 mydesign.accum\[33\] clknet_leaf_38_clk sg13g2_dfrbpq_2
XFILLER_27_701 VPWR VGND sg13g2_decap_8
XFILLER_41_214 VPWR VGND sg13g2_decap_8
XFILLER_42_759 VPWR VGND sg13g2_decap_4
XFILLER_23_973 VPWR VGND sg13g2_decap_8
XFILLER_2_811 VPWR VGND sg13g2_fill_1
X_6117__100 VPWR VGND net100 sg13g2_tiehi
XFILLER_49_314 VPWR VGND sg13g2_fill_1
XFILLER_49_303 VPWR VGND sg13g2_decap_8
XFILLER_49_347 VPWR VGND sg13g2_decap_8
XFILLER_17_200 VPWR VGND sg13g2_fill_1
XFILLER_18_756 VPWR VGND sg13g2_fill_2
XFILLER_14_984 VPWR VGND sg13g2_decap_8
X_4300_ _1240_ _1241_ _1242_ VPWR VGND sg13g2_and2_1
X_5280_ _2109_ _2094_ _2108_ VPWR VGND sg13g2_xnor2_1
X_4231_ VGND VPWR _2566_ net448 _0169_ _1179_ sg13g2_a21oi_1
XFILLER_4_52 VPWR VGND sg13g2_fill_2
XFILLER_4_63 VPWR VGND sg13g2_fill_2
X_4162_ _1106_ _1108_ _1120_ VPWR VGND sg13g2_nor2b_1
X_4093_ VGND VPWR _1058_ _1059_ _1060_ net542 sg13g2_a21oi_1
X_3113_ _2554_ net925 VPWR VGND sg13g2_inv_2
XFILLER_49_881 VPWR VGND sg13g2_decap_8
X_4995_ _1847_ _1846_ _1849_ VPWR VGND sg13g2_xor2_1
XFILLER_23_236 VPWR VGND sg13g2_decap_8
X_3946_ _0923_ _0924_ _0925_ _0926_ VPWR VGND sg13g2_or3_1
XFILLER_32_770 VPWR VGND sg13g2_fill_1
X_3877_ _0865_ _0857_ _0867_ VPWR VGND sg13g2_xor2_1
XFILLER_20_954 VPWR VGND sg13g2_decap_8
X_5616_ VGND VPWR net586 _2405_ _0327_ _2406_ sg13g2_a21oi_1
X_5547_ net481 VPWR _2347_ VGND net592 net1052 sg13g2_o21ai_1
X_5478_ mydesign.pe_weights\[22\] mydesign.pe_inputs\[9\] mydesign.accum\[11\] _2281_
+ VPWR VGND sg13g2_a21o_1
X_4429_ _1332_ _1334_ _1353_ _1355_ VPWR VGND sg13g2_or3_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
Xfanout433 net435 net433 VPWR VGND sg13g2_buf_8
Xfanout444 net445 net444 VPWR VGND sg13g2_buf_8
Xfanout466 net483 net466 VPWR VGND sg13g2_buf_8
XFILLER_24_1016 VPWR VGND sg13g2_decap_8
XFILLER_24_1027 VPWR VGND sg13g2_fill_2
Xfanout455 _0498_ net455 VPWR VGND sg13g2_buf_8
XFILLER_46_306 VPWR VGND sg13g2_fill_2
Xfanout499 _2516_ net499 VPWR VGND sg13g2_buf_8
Xfanout477 net478 net477 VPWR VGND sg13g2_buf_8
XFILLER_19_509 VPWR VGND sg13g2_fill_1
Xfanout488 net490 net488 VPWR VGND sg13g2_buf_1
X_5791__159 VPWR VGND net159 sg13g2_tiehi
XFILLER_15_759 VPWR VGND sg13g2_decap_4
XFILLER_23_781 VPWR VGND sg13g2_fill_2
XFILLER_11_954 VPWR VGND sg13g2_decap_8
XFILLER_7_936 VPWR VGND sg13g2_fill_2
X_5858__57 VPWR VGND net57 sg13g2_tiehi
XFILLER_49_122 VPWR VGND sg13g2_decap_4
X_5873__27 VPWR VGND net27 sg13g2_tiehi
X_6054__242 VPWR VGND net242 sg13g2_tiehi
XFILLER_38_807 VPWR VGND sg13g2_decap_4
XFILLER_49_177 VPWR VGND sg13g2_decap_8
XFILLER_46_873 VPWR VGND sg13g2_decap_8
XFILLER_45_394 VPWR VGND sg13g2_fill_2
X_3800_ _0796_ _0793_ _0795_ VPWR VGND sg13g2_nand2_2
X_4780_ _1658_ _1659_ _1660_ _1661_ VPWR VGND sg13g2_nor3_1
X_5926__305 VPWR VGND net305 sg13g2_tiehi
X_3731_ _0740_ _0731_ _0739_ VPWR VGND sg13g2_nand2_1
XFILLER_20_206 VPWR VGND sg13g2_fill_1
XFILLER_13_291 VPWR VGND sg13g2_fill_2
Xclkload10 clknet_leaf_21_clk clkload10/X VPWR VGND sg13g2_buf_8
X_3662_ _0674_ mydesign.accum\[114\] net540 _0653_ VPWR VGND sg13g2_and3_2
X_3593_ VGND VPWR _0512_ _0526_ _0617_ mydesign.accum\[126\] sg13g2_a21oi_1
X_5401_ _2191_ VPWR _2214_ VGND _2190_ _2193_ sg13g2_o21ai_1
X_5332_ net522 mydesign.pe_weights\[24\] net758 _2149_ VPWR VGND _2147_ sg13g2_nand4_1
XFILLER_47_1027 VPWR VGND sg13g2_fill_2
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_5263_ net464 VPWR _2093_ VGND net565 net1012 sg13g2_o21ai_1
X_4214_ _1159_ VPWR _1169_ VGND _2572_ _1157_ sg13g2_o21ai_1
X_5194_ _2027_ _2025_ _2026_ VPWR VGND sg13g2_nand2_1
X_4145_ _1101_ _1102_ _1103_ _1104_ VPWR VGND sg13g2_or3_1
X_6033__326 VPWR VGND net326 sg13g2_tiehi
X_4076_ _1043_ VPWR _1046_ VGND net543 _1045_ sg13g2_o21ai_1
XFILLER_24_512 VPWR VGND sg13g2_decap_8
XFILLER_34_49 VPWR VGND sg13g2_decap_8
X_4978_ VGND VPWR net585 _1831_ _0263_ _1832_ sg13g2_a21oi_1
Xclkload4 clknet_3_6__leaf_clk clkload4/X VPWR VGND sg13g2_buf_8
X_3929_ _2670_ net792 _0911_ _0135_ VPWR VGND sg13g2_mux2_1
XFILLER_20_762 VPWR VGND sg13g2_fill_2
X_5977__203 VPWR VGND net203 sg13g2_tiehi
XFILLER_15_501 VPWR VGND sg13g2_fill_1
XFILLER_27_350 VPWR VGND sg13g2_decap_8
XFILLER_43_865 VPWR VGND sg13g2_decap_8
XFILLER_6_298 VPWR VGND sg13g2_fill_1
XFILLER_41_7 VPWR VGND sg13g2_fill_1
XFILLER_37_125 VPWR VGND sg13g2_decap_4
XFILLER_46_670 VPWR VGND sg13g2_decap_8
X_5950_ net257 VGND VPWR _0176_ mydesign.accum\[84\] clknet_leaf_25_clk sg13g2_dfrbpq_2
XFILLER_19_873 VPWR VGND sg13g2_fill_2
X_4901_ VGND VPWR _1767_ _1769_ _0248_ net845 sg13g2_a21oi_1
XFILLER_18_372 VPWR VGND sg13g2_fill_2
XFILLER_21_504 VPWR VGND sg13g2_fill_2
X_5881_ net387 VGND VPWR _0107_ mydesign.accum\[115\] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_34_876 VPWR VGND sg13g2_fill_1
X_4832_ VGND VPWR _1710_ _1709_ _1706_ sg13g2_or2_1
XFILLER_21_537 VPWR VGND sg13g2_decap_8
XFILLER_33_386 VPWR VGND sg13g2_fill_1
X_4763_ VGND VPWR _2538_ net493 _0230_ _1650_ sg13g2_a21oi_1
XFILLER_14_1026 VPWR VGND sg13g2_fill_2
X_3714_ _0703_ _0722_ _0700_ _0724_ VPWR VGND sg13g2_nand3_1
X_4694_ _1589_ _1572_ _1588_ VPWR VGND sg13g2_nand2_1
X_3645_ VGND VPWR _2564_ net492 _0103_ _0659_ sg13g2_a21oi_1
X_3576_ _0506_ _0526_ _0601_ VPWR VGND sg13g2_and2_1
X_5315_ VGND VPWR _2527_ net449 _0296_ _2136_ sg13g2_a21oi_1
X_5246_ _2076_ _2065_ _2067_ VPWR VGND sg13g2_nand2_1
Xhold27 mydesign.inputs\[3\]\[12\] VPWR VGND net646 sg13g2_dlygate4sd3_1
Xhold16 mydesign.inputs\[3\]\[14\] VPWR VGND net422 sg13g2_dlygate4sd3_1
Xhold38 _0295_ VPWR VGND net657 sg13g2_dlygate4sd3_1
X_5177_ net459 VPWR _2013_ VGND net549 mydesign.inputs\[3\]\[10\] sg13g2_o21ai_1
Xhold49 _0015_ VPWR VGND net668 sg13g2_dlygate4sd3_1
X_4128_ _1088_ _1070_ _1086_ VPWR VGND sg13g2_xnor2_1
X_4059_ _1031_ _1015_ _1029_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_854 VPWR VGND sg13g2_fill_1
X_6109__216 VPWR VGND net216 sg13g2_tiehi
XFILLER_36_191 VPWR VGND sg13g2_fill_1
XFILLER_12_526 VPWR VGND sg13g2_decap_8
XFILLER_24_375 VPWR VGND sg13g2_fill_2
XFILLER_40_868 VPWR VGND sg13g2_decap_8
XFILLER_12_559 VPWR VGND sg13g2_fill_2
XFILLER_48_902 VPWR VGND sg13g2_decap_8
XFILLER_0_964 VPWR VGND sg13g2_decap_8
XFILLER_48_979 VPWR VGND sg13g2_decap_8
XFILLER_47_467 VPWR VGND sg13g2_fill_2
XFILLER_43_640 VPWR VGND sg13g2_decap_4
XFILLER_37_1015 VPWR VGND sg13g2_decap_8
XFILLER_43_673 VPWR VGND sg13g2_decap_8
XFILLER_15_364 VPWR VGND sg13g2_fill_1
XFILLER_31_846 VPWR VGND sg13g2_fill_2
X_3430_ net516 mydesign.accum\[54\] _0474_ VPWR VGND sg13g2_nor2b_1
X_3361_ VGND VPWR mydesign.accum\[8\] net514 _0411_ _0410_ sg13g2_a21oi_1
X_6080_ net72 VGND VPWR _0306_ mydesign.accum\[22\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_5100_ _1942_ mydesign.pe_weights\[33\] mydesign.pe_inputs\[23\] VPWR VGND sg13g2_nand2_1
X_3292_ _2688_ _2588_ _2647_ VPWR VGND sg13g2_nand2_1
X_5031_ net480 VPWR _1883_ VGND net591 net963 sg13g2_o21ai_1
XFILLER_39_935 VPWR VGND sg13g2_decap_8
XFILLER_38_412 VPWR VGND sg13g2_fill_1
Xheichips25_template_18 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_38_456 VPWR VGND sg13g2_fill_1
XFILLER_38_489 VPWR VGND sg13g2_fill_2
X_5842__85 VPWR VGND net85 sg13g2_tiehi
X_5933_ net291 VGND VPWR _0159_ mydesign.accum\[91\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_5864_ net45 VGND VPWR _0090_ mydesign.accum\[122\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_21_345 VPWR VGND sg13g2_decap_8
X_4815_ _1686_ _1693_ _1694_ VPWR VGND sg13g2_nor2_1
X_5795_ net155 VGND VPWR _0021_ mydesign.inputs\[1\]\[8\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_4746_ _1623_ _1637_ _1638_ VPWR VGND sg13g2_nor2_1
X_4677_ _1572_ _1562_ _1564_ VPWR VGND sg13g2_nand2_1
X_3628_ _0645_ mydesign.weights\[1\]\[13\] _0394_ VPWR VGND sg13g2_nand2_1
X_3559_ _0584_ _0581_ _0585_ VPWR VGND sg13g2_xor2_1
X_5229_ _2058_ _2057_ _2056_ _2060_ VPWR VGND sg13g2_a21o_1
XFILLER_29_423 VPWR VGND sg13g2_fill_1
XFILLER_29_434 VPWR VGND sg13g2_fill_1
XFILLER_45_905 VPWR VGND sg13g2_decap_8
XFILLER_16_139 VPWR VGND sg13g2_fill_2
XFILLER_40_654 VPWR VGND sg13g2_decap_8
XFILLER_9_828 VPWR VGND sg13g2_fill_2
XFILLER_48_776 VPWR VGND sg13g2_decap_8
XFILLER_47_242 VPWR VGND sg13g2_decap_4
X_6077__96 VPWR VGND net96 sg13g2_tiehi
XFILLER_36_916 VPWR VGND sg13g2_decap_8
XFILLER_44_960 VPWR VGND sg13g2_decap_8
X_4600_ net473 VPWR _1508_ VGND net574 net894 sg13g2_o21ai_1
X_5580_ VGND VPWR net587 _2371_ _0325_ _2372_ sg13g2_a21oi_1
XFILLER_7_41 VPWR VGND sg13g2_fill_1
X_4531_ _1442_ mydesign.pe_weights\[50\] mydesign.pe_inputs\[37\] VPWR VGND sg13g2_nand2_1
Xhold316 _0309_ VPWR VGND net935 sg13g2_dlygate4sd3_1
Xhold305 _0286_ VPWR VGND net924 sg13g2_dlygate4sd3_1
X_4462_ _1368_ _1384_ _1365_ _1386_ VPWR VGND sg13g2_nand3_1
X_3413_ mydesign.accum\[125\] mydesign.accum\[93\] net511 _0458_ VPWR VGND sg13g2_mux2_1
Xhold349 mydesign.accum\[101\] VPWR VGND net968 sg13g2_dlygate4sd3_1
Xhold327 mydesign.pe_inputs\[7\] VPWR VGND net946 sg13g2_dlygate4sd3_1
Xhold338 _0167_ VPWR VGND net957 sg13g2_dlygate4sd3_1
X_4393_ _1321_ _1305_ _1320_ VPWR VGND sg13g2_xnor2_1
X_3344_ _0395_ net459 _0398_ VPWR VGND sg13g2_nor2_1
X_6132_ net348 VGND VPWR _0358_ mydesign.weights\[0\]\[22\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3275_ net616 _2678_ net703 _2681_ VPWR VGND sg13g2_nand3_1
X_6063_ net206 VGND VPWR _0289_ mydesign.accum\[29\] clknet_leaf_7_clk sg13g2_dfrbpq_2
XFILLER_39_732 VPWR VGND sg13g2_fill_1
X_5014_ _1867_ _1848_ _1851_ _1866_ VPWR VGND sg13g2_and3_1
XFILLER_39_765 VPWR VGND sg13g2_decap_4
XFILLER_27_916 VPWR VGND sg13g2_fill_2
XFILLER_27_927 VPWR VGND sg13g2_decap_8
X_5934__289 VPWR VGND net289 sg13g2_tiehi
X_6083__44 VPWR VGND net44 sg13g2_tiehi
XFILLER_42_919 VPWR VGND sg13g2_decap_8
XFILLER_26_459 VPWR VGND sg13g2_decap_8
X_5916_ net325 VGND VPWR net848 mydesign.accum\[98\] clknet_leaf_44_clk sg13g2_dfrbpq_2
XFILLER_35_971 VPWR VGND sg13g2_decap_8
XFILLER_22_643 VPWR VGND sg13g2_fill_1
X_5847_ net75 VGND VPWR _0073_ net13 clknet_leaf_42_clk sg13g2_dfrbpq_2
X_5778_ net177 VGND VPWR net753 mydesign.weights\[2\]\[7\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_22_698 VPWR VGND sg13g2_decap_8
X_4729_ _1620_ _1619_ _1622_ VPWR VGND sg13g2_xor2_1
XFILLER_27_1025 VPWR VGND sg13g2_decap_4
XFILLER_29_220 VPWR VGND sg13g2_fill_2
XFILLER_45_702 VPWR VGND sg13g2_decap_8
XFILLER_44_201 VPWR VGND sg13g2_fill_1
XFILLER_17_426 VPWR VGND sg13g2_fill_1
XFILLER_29_286 VPWR VGND sg13g2_fill_1
XFILLER_45_779 VPWR VGND sg13g2_decap_8
XFILLER_26_960 VPWR VGND sg13g2_decap_8
XFILLER_41_930 VPWR VGND sg13g2_decap_8
XFILLER_40_451 VPWR VGND sg13g2_decap_4
X_5985__187 VPWR VGND net187 sg13g2_tiehi
XFILLER_12_186 VPWR VGND sg13g2_fill_2
XFILLER_48_551 VPWR VGND sg13g2_fill_1
XFILLER_36_702 VPWR VGND sg13g2_fill_1
XFILLER_17_971 VPWR VGND sg13g2_decap_8
X_3962_ VPWR _0939_ _0938_ VGND sg13g2_inv_1
X_5701_ net717 _2476_ net613 _2478_ VPWR VGND sg13g2_nand3_1
X_3893_ _0860_ VPWR _0882_ VGND _0859_ _0862_ sg13g2_o21ai_1
XFILLER_32_985 VPWR VGND sg13g2_decap_8
X_5632_ _2422_ _2408_ _2421_ VPWR VGND sg13g2_xnor2_1
X_5563_ _2359_ net650 _2356_ VPWR VGND sg13g2_nand2_1
XFILLER_8_680 VPWR VGND sg13g2_decap_8
X_4514_ net532 mydesign.pe_weights\[50\] mydesign.accum\[66\] _1426_ VPWR VGND sg13g2_a21o_1
Xhold124 _0054_ VPWR VGND net743 sg13g2_dlygate4sd3_1
Xhold113 _0343_ VPWR VGND net732 sg13g2_dlygate4sd3_1
X_5494_ _2296_ net520 mydesign.pe_weights\[21\] VPWR VGND sg13g2_nand2_1
Xhold135 mydesign.inputs\[0\]\[24\] VPWR VGND net754 sg13g2_dlygate4sd3_1
Xhold102 mydesign.accum\[120\] VPWR VGND net721 sg13g2_dlygate4sd3_1
Xhold157 mydesign.inputs\[1\]\[18\] VPWR VGND net776 sg13g2_dlygate4sd3_1
Xhold168 mydesign.inputs\[0\]\[15\] VPWR VGND net787 sg13g2_dlygate4sd3_1
X_4445_ _1347_ VPWR _1370_ VGND _1346_ _1349_ sg13g2_o21ai_1
Xhold146 mydesign.inputs\[0\]\[12\] VPWR VGND net765 sg13g2_dlygate4sd3_1
Xhold179 mydesign.inputs\[1\]\[23\] VPWR VGND net798 sg13g2_dlygate4sd3_1
X_4376_ mydesign.pe_weights\[52\] net534 net684 _1305_ VPWR VGND _1303_ sg13g2_nand4_1
Xfanout615 net619 net615 VPWR VGND sg13g2_buf_8
Xfanout604 _2625_ net604 VPWR VGND sg13g2_buf_8
X_3327_ net563 VPWR _0384_ VGND _2597_ _2598_ sg13g2_o21ai_1
X_6115_ net132 VGND VPWR net718 mydesign.weights\[3\]\[1\] clknet_leaf_49_clk sg13g2_dfrbpq_1
Xfanout637 net639 net637 VPWR VGND sg13g2_buf_8
Xfanout626 net627 net626 VPWR VGND sg13g2_buf_8
X_3258_ net769 _2668_ _2672_ _0026_ VPWR VGND sg13g2_mux2_1
X_6046_ net274 VGND VPWR net735 mydesign.accum\[32\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_2_1027 VPWR VGND sg13g2_fill_2
X_3189_ _2625_ net1 net620 VPWR VGND sg13g2_nand2_2
XFILLER_27_757 VPWR VGND sg13g2_decap_8
XFILLER_42_738 VPWR VGND sg13g2_decap_8
X_6069__188 VPWR VGND net188 sg13g2_tiehi
XFILLER_23_952 VPWR VGND sg13g2_decap_8
XFILLER_10_657 VPWR VGND sg13g2_fill_1
XFILLER_10_646 VPWR VGND sg13g2_decap_8
X_6076__104 VPWR VGND net104 sg13g2_tiehi
XFILLER_40_1022 VPWR VGND sg13g2_decap_8
XFILLER_27_93 VPWR VGND sg13g2_decap_8
XFILLER_14_963 VPWR VGND sg13g2_decap_8
X_4230_ net631 VPWR _1179_ VGND net856 net448 sg13g2_o21ai_1
X_4161_ VGND VPWR net500 _2574_ _0159_ _1119_ sg13g2_a21oi_1
X_5894__365 VPWR VGND net365 sg13g2_tiehi
XFILLER_49_860 VPWR VGND sg13g2_decap_8
X_4092_ _1059_ _0390_ mydesign.inputs\[1\]\[23\] _2595_ mydesign.inputs\[1\]\[19\]
+ VPWR VGND sg13g2_a22oi_1
X_3112_ _2553_ net537 VPWR VGND sg13g2_inv_2
XFILLER_24_727 VPWR VGND sg13g2_fill_1
X_4994_ _1848_ _1846_ _1847_ VPWR VGND sg13g2_nand2_1
X_3945_ _0925_ mydesign.weights\[3\]\[14\] net547 _0392_ VPWR VGND sg13g2_and3_1
XFILLER_17_1013 VPWR VGND sg13g2_decap_8
XFILLER_20_933 VPWR VGND sg13g2_decap_8
X_5615_ net476 VPWR _2406_ VGND net586 net1045 sg13g2_o21ai_1
X_3876_ _0857_ _0865_ _0866_ VPWR VGND sg13g2_nor2_1
X_5546_ _2346_ _2345_ _2344_ VPWR VGND sg13g2_nand2b_1
X_5477_ mydesign.pe_inputs\[9\] mydesign.pe_weights\[22\] mydesign.accum\[11\] _2280_
+ VPWR VGND sg13g2_nand3_1
X_4428_ _1353_ VPWR _1354_ VGND _1332_ _1334_ sg13g2_o21ai_1
X_4359_ VGND VPWR _2559_ net446 _0184_ _1292_ sg13g2_a21oi_1
Xfanout434 net435 net434 VPWR VGND sg13g2_buf_1
Xfanout445 net446 net445 VPWR VGND sg13g2_buf_8
Xfanout456 _0407_ net456 VPWR VGND sg13g2_buf_8
Xfanout478 net483 net478 VPWR VGND sg13g2_buf_8
Xfanout489 net490 net489 VPWR VGND sg13g2_buf_8
Xfanout467 net469 net467 VPWR VGND sg13g2_buf_8
X_6029_ net346 VGND VPWR net975 mydesign.pe_inputs\[23\] clknet_leaf_38_clk sg13g2_dfrbpq_2
XFILLER_39_381 VPWR VGND sg13g2_fill_2
XFILLER_42_546 VPWR VGND sg13g2_decap_8
XFILLER_23_771 VPWR VGND sg13g2_decap_4
XFILLER_10_443 VPWR VGND sg13g2_fill_2
XFILLER_10_454 VPWR VGND sg13g2_fill_2
XFILLER_8_0 VPWR VGND sg13g2_fill_1
XFILLER_29_9 VPWR VGND sg13g2_fill_1
XFILLER_49_189 VPWR VGND sg13g2_decap_8
XFILLER_46_852 VPWR VGND sg13g2_decap_8
XFILLER_18_543 VPWR VGND sg13g2_fill_2
XFILLER_33_502 VPWR VGND sg13g2_fill_2
XFILLER_45_373 VPWR VGND sg13g2_decap_8
X_3730_ _0739_ _0736_ _0737_ VPWR VGND sg13g2_xnor2_1
X_6061__214 VPWR VGND net214 sg13g2_tiehi
XFILLER_9_230 VPWR VGND sg13g2_decap_4
X_3661_ _0673_ mydesign.pe_inputs\[62\] _0643_ VPWR VGND sg13g2_nand2_1
X_3592_ _0512_ _0526_ mydesign.accum\[126\] _0616_ VPWR VGND sg13g2_nand3_1
X_5400_ _2211_ _2208_ _2213_ VPWR VGND sg13g2_xor2_1
Xclkload11 VPWR clkload11/Y clknet_leaf_39_clk VGND sg13g2_inv_1
X_5331_ net522 mydesign.pe_weights\[24\] net758 _2148_ VPWR VGND sg13g2_nand3_1
XFILLER_47_1006 VPWR VGND sg13g2_decap_8
X_5262_ _2092_ _2075_ _2091_ VPWR VGND sg13g2_xnor2_1
X_4213_ VGND VPWR _1164_ _1165_ _1168_ _1162_ sg13g2_a21oi_1
X_5193_ _2004_ mydesign.pe_weights\[29\] mydesign.accum\[25\] _2026_ VPWR VGND sg13g2_a21o_1
X_4144_ VGND VPWR mydesign.pe_weights\[63\] _1046_ _1103_ mydesign.accum\[91\] sg13g2_a21oi_1
X_5790__160 VPWR VGND net160 sg13g2_tiehi
X_4075_ VPWR VGND mydesign.inputs\[1\]\[20\] _1044_ net461 mydesign.inputs\[1\]\[16\]
+ _1045_ net495 sg13g2_a221oi_1
XFILLER_37_896 VPWR VGND sg13g2_decap_8
XFILLER_24_546 VPWR VGND sg13g2_decap_8
XFILLER_24_557 VPWR VGND sg13g2_fill_2
XFILLER_24_579 VPWR VGND sg13g2_fill_1
X_4977_ net474 VPWR _1832_ VGND net585 net902 sg13g2_o21ai_1
Xclkload5 clknet_3_7__leaf_clk clkload5/X VPWR VGND sg13g2_buf_8
X_3928_ _2669_ net785 _0911_ _0134_ VPWR VGND sg13g2_mux2_1
X_3859_ _0850_ _0836_ _0849_ VPWR VGND sg13g2_xnor2_1
X_5529_ VGND VPWR _2310_ _2313_ _2330_ _2328_ sg13g2_a21oi_1
XFILLER_8_1022 VPWR VGND sg13g2_decap_8
XFILLER_47_649 VPWR VGND sg13g2_decap_8
XFILLER_28_852 VPWR VGND sg13g2_fill_2
XFILLER_28_874 VPWR VGND sg13g2_fill_2
XFILLER_43_844 VPWR VGND sg13g2_decap_8
XFILLER_42_354 VPWR VGND sg13g2_decap_8
X_5839__91 VPWR VGND net91 sg13g2_tiehi
XFILLER_37_148 VPWR VGND sg13g2_decap_8
XFILLER_18_362 VPWR VGND sg13g2_fill_1
X_4900_ net612 VPWR _1770_ VGND net844 _1767_ sg13g2_o21ai_1
XFILLER_33_321 VPWR VGND sg13g2_fill_2
X_5880_ net389 VGND VPWR net878 mydesign.accum\[114\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_6008__58 VPWR VGND net58 sg13g2_tiehi
XFILLER_45_192 VPWR VGND sg13g2_decap_8
X_4831_ _1709_ _1707_ _1708_ VPWR VGND sg13g2_nand2_1
XFILLER_14_1005 VPWR VGND sg13g2_decap_8
X_4762_ net637 VPWR _1650_ VGND mydesign.pe_inputs\[30\] net493 sg13g2_o21ai_1
XFILLER_33_398 VPWR VGND sg13g2_fill_1
X_4693_ _1588_ _1573_ _1586_ VPWR VGND sg13g2_xnor2_1
X_3713_ VGND VPWR _0700_ _0703_ _0723_ _0722_ sg13g2_a21oi_1
X_3644_ net630 VPWR _0659_ VGND net492 _0658_ sg13g2_o21ai_1
X_3575_ _0600_ _0512_ _0523_ VPWR VGND sg13g2_nand2_1
X_5314_ net638 VPWR _2136_ VGND net521 net450 sg13g2_o21ai_1
X_5245_ _2070_ VPWR _2075_ VGND _2051_ _2071_ sg13g2_o21ai_1
Xhold28 mydesign.weights\[0\]\[20\] VPWR VGND net647 sg13g2_dlygate4sd3_1
Xhold17 mydesign.inputs\[2\]\[8\] VPWR VGND net423 sg13g2_dlygate4sd3_1
X_5176_ net497 mydesign.inputs\[3\]\[6\] _2012_ VPWR VGND sg13g2_nor2_1
Xhold39 mydesign.inputs\[3\]\[9\] VPWR VGND net658 sg13g2_dlygate4sd3_1
XFILLER_21_1009 VPWR VGND sg13g2_decap_8
XFILLER_28_104 VPWR VGND sg13g2_fill_1
X_4127_ _1087_ _1086_ _1070_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_126 VPWR VGND sg13g2_decap_8
X_5860__53 VPWR VGND net53 sg13g2_tiehi
X_4058_ _1030_ _1029_ _1015_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_682 VPWR VGND sg13g2_fill_1
XFILLER_12_505 VPWR VGND sg13g2_decap_8
XFILLER_20_560 VPWR VGND sg13g2_fill_2
X_5944__269 VPWR VGND net269 sg13g2_tiehi
XFILLER_20_593 VPWR VGND sg13g2_decap_8
XFILLER_0_943 VPWR VGND sg13g2_decap_8
XFILLER_48_958 VPWR VGND sg13g2_decap_8
XFILLER_31_836 VPWR VGND sg13g2_fill_1
XFILLER_35_71 VPWR VGND sg13g2_decap_4
XFILLER_31_858 VPWR VGND sg13g2_fill_2
XFILLER_7_520 VPWR VGND sg13g2_fill_1
XFILLER_7_597 VPWR VGND sg13g2_fill_1
X_3360_ net514 mydesign.accum\[40\] _0410_ VPWR VGND sg13g2_nor2b_1
XFILLER_44_1009 VPWR VGND sg13g2_decap_8
X_3291_ _2670_ net798 _2687_ _0044_ VPWR VGND sg13g2_mux2_1
X_5030_ VGND VPWR _1880_ _1881_ _1882_ net502 sg13g2_a21oi_1
XFILLER_39_914 VPWR VGND sg13g2_decap_8
Xheichips25_template_19 VPWR VGND uio_out[4] sg13g2_tielo
X_5932_ net293 VGND VPWR net965 mydesign.accum\[90\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_25_118 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_45_clk clknet_3_4__leaf_clk clknet_leaf_45_clk VPWR VGND sg13g2_buf_8
X_5863_ net47 VGND VPWR _0089_ mydesign.accum\[121\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_5794_ net156 VGND VPWR _0020_ mydesign.inputs\[2\]\[7\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_4814_ _1691_ _1670_ _1693_ VPWR VGND sg13g2_xor2_1
X_4745_ _1637_ _1621_ _1635_ VPWR VGND sg13g2_xnor2_1
X_4676_ _1566_ _1568_ _1571_ VPWR VGND sg13g2_and2_1
X_3627_ VGND VPWR _2567_ net488 _0100_ _0644_ sg13g2_a21oi_1
X_3558_ _0584_ _0582_ _0583_ VPWR VGND sg13g2_nand2_1
XFILLER_0_217 VPWR VGND sg13g2_fill_2
X_3489_ VGND VPWR _2577_ net484 _0085_ _0521_ sg13g2_a21oi_1
XFILLER_5_1014 VPWR VGND sg13g2_decap_8
X_5228_ _2057_ _2058_ _2056_ _2059_ VPWR VGND sg13g2_nand3_1
X_5159_ net474 VPWR _1998_ VGND net575 net889 sg13g2_o21ai_1
XFILLER_44_427 VPWR VGND sg13g2_fill_2
XFILLER_16_107 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_36_clk clknet_3_5__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_13_814 VPWR VGND sg13g2_decap_4
XFILLER_13_858 VPWR VGND sg13g2_fill_2
XFILLER_48_755 VPWR VGND sg13g2_decap_8
XFILLER_35_416 VPWR VGND sg13g2_decap_8
XFILLER_35_438 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_27_clk clknet_3_7__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_43_460 VPWR VGND sg13g2_fill_2
XFILLER_30_143 VPWR VGND sg13g2_fill_2
X_4530_ _1441_ mydesign.pe_weights\[49\] mydesign.pe_inputs\[38\] VPWR VGND sg13g2_nand2_1
Xhold306 mydesign.pe_weights\[50\] VPWR VGND net925 sg13g2_dlygate4sd3_1
X_4461_ VGND VPWR _1365_ _1368_ _1385_ _1384_ sg13g2_a21oi_1
Xhold317 mydesign.accum\[115\] VPWR VGND net936 sg13g2_dlygate4sd3_1
Xhold328 _0311_ VPWR VGND net947 sg13g2_dlygate4sd3_1
X_3412_ VGND VPWR _0455_ _0456_ _0072_ _0457_ sg13g2_a21oi_1
Xhold339 mydesign.accum\[122\] VPWR VGND net958 sg13g2_dlygate4sd3_1
X_4392_ _1320_ _1301_ _1318_ VPWR VGND sg13g2_xnor2_1
X_6131_ net356 VGND VPWR _0357_ mydesign.weights\[0\]\[21\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3343_ _0397_ net541 VPWR VGND net546 sg13g2_nand2b_2
X_3274_ _2680_ VPWR _0034_ VGND _2519_ _2678_ sg13g2_o21ai_1
X_6062_ net210 VGND VPWR _0288_ mydesign.accum\[28\] clknet_leaf_7_clk sg13g2_dfrbpq_2
XFILLER_23_0 VPWR VGND sg13g2_fill_2
XFILLER_39_744 VPWR VGND sg13g2_fill_1
X_5013_ _1864_ _1844_ _1866_ VPWR VGND sg13g2_xor2_1
XFILLER_38_298 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_18_clk clknet_3_3__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
XFILLER_35_950 VPWR VGND sg13g2_decap_8
X_5915_ net327 VGND VPWR net1008 mydesign.accum\[97\] clknet_leaf_44_clk sg13g2_dfrbpq_2
X_5846_ net77 VGND VPWR _0072_ net12 clknet_leaf_42_clk sg13g2_dfrbpq_2
XFILLER_22_666 VPWR VGND sg13g2_fill_2
X_5777_ net179 VGND VPWR _0003_ mydesign.weights\[2\]\[6\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_5_309 VPWR VGND sg13g2_fill_2
X_4728_ _1621_ _1619_ _1620_ VPWR VGND sg13g2_nand2_1
X_4659_ _1555_ mydesign.pe_weights\[44\] _1531_ VPWR VGND sg13g2_nand2b_1
XFILLER_1_504 VPWR VGND sg13g2_fill_2
XFILLER_27_1004 VPWR VGND sg13g2_decap_8
XFILLER_18_939 VPWR VGND sg13g2_decap_8
XFILLER_45_758 VPWR VGND sg13g2_decap_8
XFILLER_44_224 VPWR VGND sg13g2_fill_1
XFILLER_41_986 VPWR VGND sg13g2_decap_8
XFILLER_40_463 VPWR VGND sg13g2_decap_8
XFILLER_34_1019 VPWR VGND sg13g2_decap_8
XFILLER_5_854 VPWR VGND sg13g2_fill_1
XFILLER_5_887 VPWR VGND sg13g2_fill_1
XFILLER_5_876 VPWR VGND sg13g2_decap_8
XFILLER_4_364 VPWR VGND sg13g2_fill_2
X_6057__230 VPWR VGND net230 sg13g2_tiehi
XFILLER_0_581 VPWR VGND sg13g2_decap_8
XFILLER_17_950 VPWR VGND sg13g2_decap_8
X_3961_ mydesign.pe_inputs\[52\] _0919_ mydesign.accum\[97\] _0938_ VPWR VGND sg13g2_nand3_1
XFILLER_35_257 VPWR VGND sg13g2_fill_1
X_5700_ _2477_ VPWR _0340_ VGND net603 _2476_ sg13g2_o21ai_1
X_3892_ _0879_ _0877_ _0881_ VPWR VGND sg13g2_xor2_1
XFILLER_32_964 VPWR VGND sg13g2_decap_8
X_5631_ _2418_ _2409_ _2421_ VPWR VGND sg13g2_xor2_1
XFILLER_31_463 VPWR VGND sg13g2_decap_8
X_5562_ _2358_ VPWR _0321_ VGND net601 _2355_ sg13g2_o21ai_1
X_4513_ mydesign.pe_weights\[50\] net532 mydesign.accum\[66\] _1425_ VPWR VGND sg13g2_nand3_1
Xhold125 mydesign.cp2\[0\] VPWR VGND net744 sg13g2_dlygate4sd3_1
Xhold114 mydesign.weights\[2\]\[5\] VPWR VGND net733 sg13g2_dlygate4sd3_1
X_5493_ VGND VPWR net588 _2294_ _0315_ _2295_ sg13g2_a21oi_1
Xhold103 mydesign.weights\[0\]\[23\] VPWR VGND net722 sg13g2_dlygate4sd3_1
Xhold147 mydesign.inputs\[0\]\[17\] VPWR VGND net766 sg13g2_dlygate4sd3_1
Xhold136 mydesign.out\[0\] VPWR VGND net755 sg13g2_dlygate4sd3_1
X_4444_ _1367_ _1364_ _1369_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_7_clk clknet_3_6__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xhold158 mydesign.weights\[1\]\[11\] VPWR VGND net777 sg13g2_dlygate4sd3_1
Xhold169 mydesign.inputs\[0\]\[18\] VPWR VGND net788 sg13g2_dlygate4sd3_1
Xfanout605 _2617_ net605 VPWR VGND sg13g2_buf_8
X_4375_ mydesign.pe_weights\[52\] net534 net684 _1304_ VPWR VGND sg13g2_nand3_1
X_6036__314 VPWR VGND net314 sg13g2_tiehi
X_3326_ net607 _0383_ _0060_ VPWR VGND sg13g2_nor2_1
X_6114_ net140 VGND VPWR net726 mydesign.weights\[3\]\[0\] clknet_leaf_49_clk sg13g2_dfrbpq_1
Xfanout616 net617 net616 VPWR VGND sg13g2_buf_8
Xfanout627 net640 net627 VPWR VGND sg13g2_buf_8
Xfanout638 net639 net638 VPWR VGND sg13g2_buf_8
X_6045_ net278 VGND VPWR net817 mydesign.pe_weights\[19\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3257_ net762 _2667_ _2672_ _0025_ VPWR VGND sg13g2_mux2_1
XFILLER_2_1006 VPWR VGND sg13g2_decap_8
X_3188_ net754 _2623_ net620 _2624_ VPWR VGND sg13g2_nand3_1
XFILLER_22_441 VPWR VGND sg13g2_fill_2
X_5829_ net111 VGND VPWR net713 mydesign.inputs\[3\]\[2\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_5_128 VPWR VGND sg13g2_fill_2
XFILLER_2_879 VPWR VGND sg13g2_fill_1
XFILLER_49_327 VPWR VGND sg13g2_decap_8
XFILLER_40_1001 VPWR VGND sg13g2_decap_8
XFILLER_18_758 VPWR VGND sg13g2_fill_1
XFILLER_14_942 VPWR VGND sg13g2_decap_8
XFILLER_43_93 VPWR VGND sg13g2_fill_2
XFILLER_40_271 VPWR VGND sg13g2_decap_4
XFILLER_13_496 VPWR VGND sg13g2_decap_8
X_4160_ net469 VPWR _1119_ VGND net499 _1118_ sg13g2_o21ai_1
XFILLER_4_65 VPWR VGND sg13g2_fill_1
X_3111_ VPWR _2552_ net815 VGND sg13g2_inv_1
X_4091_ _1058_ mydesign.inputs\[1\]\[15\] _0394_ VPWR VGND sg13g2_nand2_1
XFILLER_36_500 VPWR VGND sg13g2_fill_1
XFILLER_48_393 VPWR VGND sg13g2_fill_1
XFILLER_17_780 VPWR VGND sg13g2_decap_8
X_4993_ _1825_ VPWR _1847_ VGND _1814_ _1826_ sg13g2_o21ai_1
XFILLER_24_739 VPWR VGND sg13g2_fill_2
X_3944_ _0924_ net541 mydesign.weights\[3\]\[2\] net496 VPWR VGND sg13g2_and3_1
X_3875_ _0865_ _0858_ _0863_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_912 VPWR VGND sg13g2_decap_8
X_5614_ _2403_ _2384_ _2405_ VPWR VGND sg13g2_xor2_1
XFILLER_31_282 VPWR VGND sg13g2_fill_1
XFILLER_20_989 VPWR VGND sg13g2_decap_8
X_5545_ _2343_ VPWR _2345_ VGND _2327_ _2330_ sg13g2_o21ai_1
X_5476_ _2279_ net521 mydesign.pe_weights\[23\] VPWR VGND sg13g2_nand2_1
X_4427_ _1352_ _1344_ _1353_ VPWR VGND sg13g2_xor2_1
X_4358_ net633 VPWR _1292_ VGND net943 net446 sg13g2_o21ai_1
Xfanout446 net453 net446 VPWR VGND sg13g2_buf_8
Xfanout435 net439 net435 VPWR VGND sg13g2_buf_1
Xfanout457 net458 net457 VPWR VGND sg13g2_buf_8
X_4289_ _1214_ VPWR _1231_ VGND _1213_ _1216_ sg13g2_o21ai_1
Xfanout468 net469 net468 VPWR VGND sg13g2_buf_8
X_3309_ net712 net429 net618 _2695_ VPWR VGND sg13g2_nand3_1
Xfanout479 net480 net479 VPWR VGND sg13g2_buf_8
XFILLER_46_308 VPWR VGND sg13g2_fill_1
X_6028_ net350 VGND VPWR _0254_ mydesign.pe_inputs\[22\] clknet_leaf_38_clk sg13g2_dfrbpq_2
XFILLER_15_717 VPWR VGND sg13g2_fill_2
XFILLER_7_905 VPWR VGND sg13g2_fill_1
XFILLER_13_30 VPWR VGND sg13g2_fill_1
XFILLER_7_938 VPWR VGND sg13g2_fill_1
XFILLER_7_927 VPWR VGND sg13g2_fill_1
XFILLER_6_404 VPWR VGND sg13g2_decap_4
XFILLER_11_989 VPWR VGND sg13g2_decap_8
XFILLER_1_153 VPWR VGND sg13g2_fill_2
X_5954__249 VPWR VGND net249 sg13g2_tiehi
XFILLER_18_500 VPWR VGND sg13g2_fill_2
XFILLER_37_308 VPWR VGND sg13g2_fill_2
XFILLER_46_831 VPWR VGND sg13g2_decap_8
XFILLER_18_588 VPWR VGND sg13g2_fill_2
XFILLER_33_514 VPWR VGND sg13g2_fill_1
XFILLER_33_525 VPWR VGND sg13g2_fill_2
XFILLER_41_591 VPWR VGND sg13g2_fill_1
XFILLER_9_220 VPWR VGND sg13g2_fill_1
XFILLER_13_293 VPWR VGND sg13g2_fill_1
X_3660_ VGND VPWR net578 _0671_ _0105_ _0672_ sg13g2_a21oi_1
X_3591_ VGND VPWR mydesign.accum\[125\] _0601_ _0615_ _0603_ sg13g2_a21oi_1
Xclkload12 VPWR clkload12/Y clknet_leaf_41_clk VGND sg13g2_inv_1
X_5330_ _2145_ _2146_ _2147_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_993 VPWR VGND sg13g2_decap_8
XFILLER_5_481 VPWR VGND sg13g2_fill_2
X_5261_ _2091_ _2076_ _2089_ VPWR VGND sg13g2_xnor2_1
X_4212_ VGND VPWR net569 _1166_ _0162_ _1167_ sg13g2_a21oi_1
X_5192_ mydesign.pe_weights\[29\] _2004_ mydesign.accum\[25\] _2025_ VPWR VGND sg13g2_nand3_1
X_4143_ _1102_ mydesign.accum\[91\] mydesign.pe_weights\[63\] _1046_ VPWR VGND sg13g2_and3_1
X_4074_ _1044_ net544 net555 mydesign.inputs\[1\]\[12\] VPWR VGND sg13g2_and3_1
XFILLER_36_396 VPWR VGND sg13g2_fill_1
X_4976_ _1829_ _1812_ _1831_ VPWR VGND sg13g2_xor2_1
X_3927_ _2668_ net768 _0911_ _0133_ VPWR VGND sg13g2_mux2_1
Xclkload6 clkload6/Y clknet_leaf_49_clk VPWR VGND sg13g2_inv_2
X_3858_ _0846_ _0823_ _0849_ VPWR VGND sg13g2_xor2_1
X_3789_ net459 VPWR _0786_ VGND net550 mydesign.weights\[2\]\[9\] sg13g2_o21ai_1
XFILLER_30_1011 VPWR VGND sg13g2_decap_8
X_5528_ _2329_ _2310_ _2313_ _2328_ VPWR VGND sg13g2_and3_1
X_5459_ net525 mydesign.pe_inputs\[8\] mydesign.accum\[10\] _2263_ VPWR VGND sg13g2_a21o_1
XFILLER_8_1001 VPWR VGND sg13g2_decap_8
XFILLER_47_628 VPWR VGND sg13g2_decap_8
XFILLER_46_105 VPWR VGND sg13g2_fill_2
XFILLER_27_341 VPWR VGND sg13g2_decap_4
XFILLER_28_886 VPWR VGND sg13g2_decap_8
XFILLER_43_823 VPWR VGND sg13g2_decap_8
XFILLER_42_388 VPWR VGND sg13g2_decap_4
XFILLER_3_985 VPWR VGND sg13g2_decap_8
XFILLER_38_628 VPWR VGND sg13g2_decap_8
XFILLER_38_617 VPWR VGND sg13g2_fill_1
XFILLER_19_875 VPWR VGND sg13g2_fill_1
XFILLER_18_374 VPWR VGND sg13g2_fill_1
XFILLER_34_823 VPWR VGND sg13g2_fill_2
X_4830_ mydesign.pe_inputs\[29\] net533 mydesign.accum\[52\] _1708_ VPWR VGND sg13g2_a21o_1
XFILLER_33_344 VPWR VGND sg13g2_fill_2
XFILLER_21_506 VPWR VGND sg13g2_fill_1
X_4761_ VGND VPWR _2546_ net447 _0229_ _1649_ sg13g2_a21oi_1
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
X_4692_ _1587_ _1586_ _1573_ VPWR VGND sg13g2_nand2b_1
X_3712_ _0720_ _0710_ _0722_ VPWR VGND sg13g2_xor2_1
X_3643_ _0655_ VPWR _0658_ VGND net542 _0657_ sg13g2_o21ai_1
X_3574_ _0586_ VPWR _0599_ VGND _0579_ _0587_ sg13g2_o21ai_1
X_5313_ _2135_ VPWR _0295_ VGND net597 _2130_ sg13g2_o21ai_1
X_5244_ VGND VPWR net499 _2528_ _0287_ _2074_ sg13g2_a21oi_1
Xhold29 mydesign.inputs\[3\]\[7\] VPWR VGND net648 sg13g2_dlygate4sd3_1
X_5175_ VGND VPWR net445 _2009_ _0281_ _2011_ sg13g2_a21oi_1
Xhold18 _0013_ VPWR VGND net424 sg13g2_dlygate4sd3_1
X_4126_ _1084_ _1085_ _1086_ VPWR VGND sg13g2_nor2b_1
X_4057_ _1029_ _1026_ _1027_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_867 VPWR VGND sg13g2_fill_2
X_4959_ _1814_ mydesign.pe_weights\[36\] mydesign.pe_inputs\[27\] VPWR VGND sg13g2_nand2_1
XFILLER_0_922 VPWR VGND sg13g2_decap_8
XFILLER_48_937 VPWR VGND sg13g2_decap_8
XFILLER_0_999 VPWR VGND sg13g2_decap_8
XFILLER_47_425 VPWR VGND sg13g2_decap_4
XFILLER_47_469 VPWR VGND sg13g2_fill_1
XFILLER_16_812 VPWR VGND sg13g2_decap_4
XFILLER_28_683 VPWR VGND sg13g2_decap_4
XFILLER_15_322 VPWR VGND sg13g2_fill_1
XFILLER_27_193 VPWR VGND sg13g2_fill_2
XFILLER_42_152 VPWR VGND sg13g2_fill_1
XFILLER_31_815 VPWR VGND sg13g2_fill_2
XFILLER_31_848 VPWR VGND sg13g2_fill_1
XFILLER_7_510 VPWR VGND sg13g2_fill_1
X_3290_ _2669_ net793 _2687_ _0043_ VPWR VGND sg13g2_mux2_1
XFILLER_20_1010 VPWR VGND sg13g2_decap_8
XFILLER_47_992 VPWR VGND sg13g2_decap_8
X_5931_ net295 VGND VPWR net897 mydesign.accum\[89\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_5862_ net49 VGND VPWR _0088_ mydesign.accum\[120\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_5793_ net157 VGND VPWR _0019_ mydesign.inputs\[2\]\[6\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_4813_ _1670_ _1691_ _1692_ VPWR VGND sg13g2_nor2b_1
X_4744_ _1621_ _1635_ _1636_ VPWR VGND sg13g2_nor2_1
XFILLER_30_892 VPWR VGND sg13g2_decap_8
X_4675_ VGND VPWR net560 _1569_ _0222_ _1570_ sg13g2_a21oi_1
X_3626_ net626 VPWR _0644_ VGND net487 _0643_ sg13g2_o21ai_1
X_3557_ _0526_ _0501_ mydesign.accum\[124\] _0583_ VPWR VGND sg13g2_a21o_1
X_3488_ net621 VPWR _0521_ VGND net485 _0520_ sg13g2_o21ai_1
X_5227_ _2004_ mydesign.pe_weights\[31\] mydesign.accum\[27\] _2058_ VPWR VGND sg13g2_a21o_1
XFILLER_29_403 VPWR VGND sg13g2_decap_8
X_5158_ _1997_ _1993_ _1996_ VPWR VGND sg13g2_xnor2_1
X_4109_ mydesign.pe_weights\[61\] _1046_ mydesign.accum\[89\] _1070_ VPWR VGND sg13g2_nand3_1
X_5089_ _1924_ _1931_ _1932_ VPWR VGND sg13g2_nor2_1
XFILLER_25_653 VPWR VGND sg13g2_fill_2
XFILLER_12_314 VPWR VGND sg13g2_fill_1
XFILLER_21_96 VPWR VGND sg13g2_fill_2
XFILLER_48_734 VPWR VGND sg13g2_decap_8
XFILLER_0_796 VPWR VGND sg13g2_decap_8
XFILLER_16_642 VPWR VGND sg13g2_fill_1
XFILLER_44_995 VPWR VGND sg13g2_decap_8
XFILLER_43_472 VPWR VGND sg13g2_fill_1
XFILLER_7_351 VPWR VGND sg13g2_fill_2
XFILLER_11_380 VPWR VGND sg13g2_decap_8
Xhold307 mydesign.accum\[52\] VPWR VGND net926 sg13g2_dlygate4sd3_1
X_4460_ _1384_ _1382_ _1383_ VPWR VGND sg13g2_nand2_1
Xhold329 mydesign.accum\[95\] VPWR VGND net948 sg13g2_dlygate4sd3_1
X_4391_ _1319_ _1301_ _1318_ VPWR VGND sg13g2_nand2_1
X_3411_ net622 VPWR _0457_ VGND net1075 net430 sg13g2_o21ai_1
Xhold318 mydesign.accum\[121\] VPWR VGND net937 sg13g2_dlygate4sd3_1
X_6130_ net364 VGND VPWR _0356_ mydesign.weights\[0\]\[20\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3342_ net545 net543 _0396_ VPWR VGND sg13g2_nor2b_2
X_3273_ net617 _2678_ net682 _2680_ VPWR VGND sg13g2_nand3_1
X_6061_ net214 VGND VPWR _0287_ mydesign.accum\[27\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5012_ _1844_ _1864_ _1865_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_200 VPWR VGND sg13g2_fill_2
X_5914_ net329 VGND VPWR _0140_ mydesign.accum\[96\] clknet_leaf_44_clk sg13g2_dfrbpq_2
X_5845_ net79 VGND VPWR _0071_ net11 clknet_leaf_42_clk sg13g2_dfrbpq_2
XFILLER_22_634 VPWR VGND sg13g2_fill_1
X_5776_ net181 VGND VPWR _0002_ mydesign.weights\[2\]\[5\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_4727_ _1598_ VPWR _1620_ VGND _1597_ _1600_ sg13g2_o21ai_1
X_4658_ VGND VPWR net560 _1553_ _0221_ _1554_ sg13g2_a21oi_1
X_3609_ _0632_ _0621_ _0631_ VPWR VGND sg13g2_xnor2_1
X_4589_ net537 mydesign.pe_inputs\[39\] mydesign.accum\[70\] _1497_ VPWR VGND sg13g2_nand3_1
XFILLER_29_222 VPWR VGND sg13g2_fill_1
XFILLER_29_233 VPWR VGND sg13g2_fill_1
XFILLER_45_737 VPWR VGND sg13g2_decap_8
XFILLER_44_214 VPWR VGND sg13g2_fill_2
XFILLER_13_634 VPWR VGND sg13g2_fill_1
XFILLER_26_995 VPWR VGND sg13g2_decap_8
XFILLER_41_965 VPWR VGND sg13g2_decap_8
XFILLER_12_122 VPWR VGND sg13g2_decap_8
XFILLER_12_133 VPWR VGND sg13g2_fill_2
XFILLER_5_833 VPWR VGND sg13g2_fill_2
XFILLER_32_84 VPWR VGND sg13g2_fill_2
X_5933__291 VPWR VGND net291 sg13g2_tiehi
XFILLER_35_214 VPWR VGND sg13g2_fill_1
X_3960_ net462 net1054 _0140_ VPWR VGND sg13g2_nor2_1
XFILLER_44_792 VPWR VGND sg13g2_decap_8
XFILLER_16_472 VPWR VGND sg13g2_decap_4
XFILLER_32_943 VPWR VGND sg13g2_decap_8
X_6064__202 VPWR VGND net202 sg13g2_tiehi
X_5964__229 VPWR VGND net229 sg13g2_tiehi
X_3891_ _0877_ _0879_ _0880_ VPWR VGND sg13g2_nor2_1
X_5630_ _2409_ _2418_ _2420_ VPWR VGND sg13g2_nor2_1
X_5561_ _2358_ net658 _2356_ VPWR VGND sg13g2_nand2_1
X_4512_ _1424_ mydesign.pe_weights\[49\] mydesign.pe_inputs\[37\] VPWR VGND sg13g2_nand2_1
X_5492_ net478 VPWR _2295_ VGND net588 net970 sg13g2_o21ai_1
Xhold115 mydesign.accum\[32\] VPWR VGND net734 sg13g2_dlygate4sd3_1
Xhold104 mydesign.weights\[0\]\[24\] VPWR VGND net723 sg13g2_dlygate4sd3_1
Xhold126 mydesign.accum\[48\] VPWR VGND net745 sg13g2_dlygate4sd3_1
Xhold159 mydesign.inputs\[1\]\[19\] VPWR VGND net778 sg13g2_dlygate4sd3_1
Xhold137 mydesign.cp2\[1\] VPWR VGND net756 sg13g2_dlygate4sd3_1
X_4443_ VGND VPWR _1368_ _1367_ _1364_ sg13g2_or2_1
Xhold148 mydesign.weights\[0\]\[12\] VPWR VGND net767 sg13g2_dlygate4sd3_1
Xfanout606 _2617_ net606 VPWR VGND sg13g2_buf_8
X_4374_ _1301_ _1302_ _1303_ VPWR VGND sg13g2_nor2b_1
X_3325_ _0383_ _0380_ net1064 _2658_ _2600_ VPWR VGND sg13g2_a22oi_1
Xfanout617 net619 net617 VPWR VGND sg13g2_buf_8
Xfanout628 net632 net628 VPWR VGND sg13g2_buf_8
X_6113_ net176 VGND VPWR net1104 mydesign.out\[3\] clknet_leaf_43_clk sg13g2_dfrbpq_1
Xfanout639 net640 net639 VPWR VGND sg13g2_buf_8
X_6044_ net282 VGND VPWR _0270_ mydesign.pe_weights\[18\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3256_ net614 VPWR _2672_ VGND _2618_ _2671_ sg13g2_o21ai_1
X_3187_ _2619_ _2621_ net605 _2623_ VPWR VGND sg13g2_nand3_1
XFILLER_41_228 VPWR VGND sg13g2_fill_1
XFILLER_35_781 VPWR VGND sg13g2_decap_4
X_5828_ net113 VGND VPWR net743 mydesign.inputs\[3\]\[1\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_23_987 VPWR VGND sg13g2_decap_8
X_5759_ VGND VPWR _1775_ _2505_ _0367_ net870 sg13g2_a21oi_1
XFILLER_33_718 VPWR VGND sg13g2_fill_2
XFILLER_13_453 VPWR VGND sg13g2_fill_1
XFILLER_13_464 VPWR VGND sg13g2_fill_1
XFILLER_14_998 VPWR VGND sg13g2_decap_8
XFILLER_4_151 VPWR VGND sg13g2_decap_8
XFILLER_4_184 VPWR VGND sg13g2_decap_4
XFILLER_4_173 VPWR VGND sg13g2_fill_2
XFILLER_1_880 VPWR VGND sg13g2_decap_8
X_3110_ VPWR _2551_ net811 VGND sg13g2_inv_1
X_4090_ VGND VPWR _2569_ net489 _0150_ _1057_ sg13g2_a21oi_1
XFILLER_49_895 VPWR VGND sg13g2_decap_8
XFILLER_24_707 VPWR VGND sg13g2_decap_4
X_4992_ _1844_ _1845_ _1846_ VPWR VGND sg13g2_and2_1
X_3943_ VGND VPWR _0921_ _0922_ _0923_ _0397_ sg13g2_a21oi_1
X_6068__190 VPWR VGND net190 sg13g2_tiehi
X_3874_ _0858_ _0863_ _0864_ VPWR VGND sg13g2_and2_1
XFILLER_32_784 VPWR VGND sg13g2_fill_2
X_5613_ _2404_ _2403_ _2384_ VPWR VGND sg13g2_nand2b_1
XFILLER_20_968 VPWR VGND sg13g2_decap_8
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
X_5784__169 VPWR VGND net169 sg13g2_tiehi
XFILLER_8_490 VPWR VGND sg13g2_fill_2
XFILLER_9_991 VPWR VGND sg13g2_decap_8
X_5544_ _2327_ _2330_ _2343_ _2344_ VPWR VGND sg13g2_nor3_1
X_5475_ _2278_ mydesign.pe_inputs\[10\] mydesign.pe_weights\[21\] VPWR VGND sg13g2_nand2_1
X_4426_ _1352_ _1345_ _1350_ VPWR VGND sg13g2_xnor2_1
XFILLER_48_28 VPWR VGND sg13g2_decap_4
Xfanout436 net437 net436 VPWR VGND sg13g2_buf_8
X_4357_ VGND VPWR _2560_ net434 _0183_ _1291_ sg13g2_a21oi_1
Xfanout447 net452 net447 VPWR VGND sg13g2_buf_8
X_4288_ _1230_ mydesign.pe_weights\[57\] mydesign.pe_inputs\[47\] VPWR VGND sg13g2_nand2_1
Xfanout469 net483 net469 VPWR VGND sg13g2_buf_8
X_3308_ _2694_ VPWR _0054_ VGND net601 net429 sg13g2_o21ai_1
Xfanout458 _0403_ net458 VPWR VGND sg13g2_buf_8
X_3239_ _2658_ net605 net607 _2659_ VPWR VGND sg13g2_a21o_2
X_6027_ net354 VGND VPWR net850 mydesign.pe_inputs\[21\] clknet_leaf_35_clk sg13g2_dfrbpq_2
XFILLER_39_372 VPWR VGND sg13g2_decap_4
XFILLER_15_707 VPWR VGND sg13g2_fill_1
XFILLER_11_968 VPWR VGND sg13g2_decap_8
XFILLER_10_456 VPWR VGND sg13g2_fill_1
XFILLER_13_53 VPWR VGND sg13g2_fill_2
XFILLER_13_97 VPWR VGND sg13g2_fill_1
XFILLER_2_622 VPWR VGND sg13g2_decap_4
Xhold490 _2639_ VPWR VGND net1109 sg13g2_dlygate4sd3_1
XFILLER_49_114 VPWR VGND sg13g2_decap_4
XFILLER_49_103 VPWR VGND sg13g2_fill_2
XFILLER_49_147 VPWR VGND sg13g2_decap_8
XFILLER_49_158 VPWR VGND sg13g2_fill_1
XFILLER_46_810 VPWR VGND sg13g2_decap_8
XFILLER_46_887 VPWR VGND sg13g2_decap_8
XFILLER_45_353 VPWR VGND sg13g2_decap_4
XFILLER_18_545 VPWR VGND sg13g2_fill_1
XFILLER_33_504 VPWR VGND sg13g2_fill_1
XFILLER_14_740 VPWR VGND sg13g2_fill_1
X_6026__358 VPWR VGND net358 sg13g2_tiehi
X_3590_ VGND VPWR net558 _0613_ _0093_ _0614_ sg13g2_a21oi_1
Xclkload13 clkload13/Y clknet_leaf_32_clk VPWR VGND sg13g2_inv_2
XFILLER_6_972 VPWR VGND sg13g2_decap_8
X_5260_ VGND VPWR _2065_ _2067_ _2090_ _2089_ sg13g2_a21oi_1
X_4211_ net471 VPWR _1167_ VGND net569 net806 sg13g2_o21ai_1
X_5191_ net462 _2024_ _0284_ VPWR VGND sg13g2_nor2_1
X_4142_ _1101_ mydesign.pe_weights\[62\] _1051_ VPWR VGND sg13g2_nand2_1
XFILLER_28_309 VPWR VGND sg13g2_decap_4
X_4073_ mydesign.inputs\[1\]\[8\] net460 net498 _1043_ VPWR VGND sg13g2_nand3_1
XFILLER_49_692 VPWR VGND sg13g2_decap_8
XFILLER_37_876 VPWR VGND sg13g2_decap_4
X_4975_ _1829_ _1812_ _1830_ VPWR VGND sg13g2_nor2b_1
X_3926_ _2667_ net783 _0911_ _0132_ VPWR VGND sg13g2_mux2_1
Xclkload7 clknet_leaf_2_clk clkload7/X VPWR VGND sg13g2_buf_8
X_3857_ _0823_ _0846_ _0848_ VPWR VGND sg13g2_nor2_1
X_3788_ net497 mydesign.weights\[2\]\[5\] _0785_ VPWR VGND sg13g2_nor2_1
XFILLER_4_909 VPWR VGND sg13g2_decap_4
X_5527_ _2326_ _2306_ _2328_ VPWR VGND sg13g2_xor2_1
X_5458_ mydesign.pe_inputs\[8\] net525 mydesign.accum\[10\] _2262_ VPWR VGND sg13g2_nand3_1
X_5389_ _2201_ _2200_ _2203_ VPWR VGND sg13g2_xor2_1
X_4409_ _1336_ _1313_ _1335_ VPWR VGND sg13g2_nand2_1
X_5877__395 VPWR VGND net395 sg13g2_tiehi
XFILLER_47_607 VPWR VGND sg13g2_decap_8
XFILLER_43_802 VPWR VGND sg13g2_decap_8
XFILLER_27_364 VPWR VGND sg13g2_decap_8
XFILLER_27_386 VPWR VGND sg13g2_fill_2
XFILLER_43_879 VPWR VGND sg13g2_decap_8
XFILLER_15_559 VPWR VGND sg13g2_fill_2
XFILLER_3_964 VPWR VGND sg13g2_decap_8
XFILLER_38_607 VPWR VGND sg13g2_decap_4
XFILLER_37_139 VPWR VGND sg13g2_decap_4
XFILLER_46_684 VPWR VGND sg13g2_decap_8
XFILLER_33_301 VPWR VGND sg13g2_fill_1
XFILLER_18_397 VPWR VGND sg13g2_decap_4
X_4760_ net637 VPWR _1649_ VGND net849 net447 sg13g2_o21ai_1
X_3711_ _0721_ _0720_ VPWR VGND _0710_ sg13g2_nand2b_2
X_4691_ _1584_ _1560_ _1586_ VPWR VGND sg13g2_xor2_1
X_3642_ VPWR VGND mydesign.weights\[1\]\[23\] _0656_ net461 mydesign.weights\[1\]\[19\]
+ _0657_ net495 sg13g2_a221oi_1
X_3573_ _0598_ _0592_ _0595_ VPWR VGND sg13g2_nand2_1
X_5312_ _2135_ net656 _2131_ VPWR VGND sg13g2_nand2_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
X_5243_ net466 VPWR _2074_ VGND net499 _2073_ sg13g2_o21ai_1
X_5174_ net634 VPWR _2011_ VGND net976 net445 sg13g2_o21ai_1
Xhold19 mydesign.inputs\[2\]\[13\] VPWR VGND net425 sg13g2_dlygate4sd3_1
X_4125_ _1083_ VPWR _1085_ VGND _1081_ _1082_ sg13g2_o21ai_1
XFILLER_37_651 VPWR VGND sg13g2_fill_2
X_4056_ VPWR _1028_ _1027_ VGND sg13g2_inv_1
XFILLER_25_879 VPWR VGND sg13g2_decap_4
X_4958_ _1804_ VPWR _1813_ VGND _1797_ _1805_ sg13g2_o21ai_1
X_4889_ _1763_ net654 _1762_ VPWR VGND sg13g2_nand2_1
X_3909_ _0897_ _0895_ _0896_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_901 VPWR VGND sg13g2_decap_8
XFILLER_48_916 VPWR VGND sg13g2_decap_8
XFILLER_0_978 VPWR VGND sg13g2_decap_8
XFILLER_15_345 VPWR VGND sg13g2_fill_2
XFILLER_16_857 VPWR VGND sg13g2_fill_2
XFILLER_43_687 VPWR VGND sg13g2_decap_8
XFILLER_42_131 VPWR VGND sg13g2_decap_4
XFILLER_15_378 VPWR VGND sg13g2_decap_8
XFILLER_30_304 VPWR VGND sg13g2_decap_8
XFILLER_24_890 VPWR VGND sg13g2_fill_2
XFILLER_30_315 VPWR VGND sg13g2_fill_1
XFILLER_11_540 VPWR VGND sg13g2_fill_1
XFILLER_30_348 VPWR VGND sg13g2_fill_2
X_5995__114 VPWR VGND net114 sg13g2_tiehi
XFILLER_39_949 VPWR VGND sg13g2_decap_8
XFILLER_38_437 VPWR VGND sg13g2_fill_2
XFILLER_19_651 VPWR VGND sg13g2_fill_1
XFILLER_47_971 VPWR VGND sg13g2_decap_8
X_5930_ net297 VGND VPWR _0156_ mydesign.accum\[88\] clknet_leaf_16_clk sg13g2_dfrbpq_2
XFILLER_46_481 VPWR VGND sg13g2_fill_1
X_5861_ net51 VGND VPWR _0087_ mydesign.pe_weights\[63\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_22_805 VPWR VGND sg13g2_fill_2
X_5792_ net158 VGND VPWR _0018_ mydesign.inputs\[2\]\[5\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_33_175 VPWR VGND sg13g2_fill_1
X_4812_ _1690_ _1687_ _1691_ VPWR VGND sg13g2_xor2_1
XFILLER_21_359 VPWR VGND sg13g2_decap_4
X_4743_ _1635_ _1633_ _1634_ VPWR VGND sg13g2_xnor2_1
X_5943__271 VPWR VGND net271 sg13g2_tiehi
X_4674_ net467 VPWR _1570_ VGND net560 net959 sg13g2_o21ai_1
X_3625_ _0639_ net802 _0642_ _0643_ VPWR VGND sg13g2_a21o_2
X_3556_ _0501_ _0526_ mydesign.accum\[124\] _0582_ VPWR VGND sg13g2_nand3_1
XFILLER_1_709 VPWR VGND sg13g2_fill_1
X_6039__302 VPWR VGND net302 sg13g2_tiehi
X_5974__209 VPWR VGND net209 sg13g2_tiehi
X_5226_ mydesign.pe_weights\[31\] _2004_ mydesign.accum\[27\] _2057_ VPWR VGND sg13g2_nand3_1
X_3487_ _2586_ _0519_ _0520_ VPWR VGND sg13g2_and2_1
X_5157_ _1996_ _1994_ _1995_ VPWR VGND sg13g2_xnor2_1
X_4108_ net462 _1069_ _0156_ VPWR VGND sg13g2_nor2_1
XFILLER_45_919 VPWR VGND sg13g2_decap_8
X_5088_ _1929_ _1908_ _1931_ VPWR VGND sg13g2_xor2_1
XFILLER_44_429 VPWR VGND sg13g2_fill_1
XFILLER_38_993 VPWR VGND sg13g2_decap_8
X_4039_ _1012_ _1010_ _1011_ VPWR VGND sg13g2_nand2_1
XFILLER_25_676 VPWR VGND sg13g2_fill_2
XFILLER_40_668 VPWR VGND sg13g2_decap_8
XFILLER_12_337 VPWR VGND sg13g2_decap_4
XFILLER_4_503 VPWR VGND sg13g2_decap_8
XFILLER_48_713 VPWR VGND sg13g2_decap_8
XFILLER_0_775 VPWR VGND sg13g2_decap_8
XFILLER_29_993 VPWR VGND sg13g2_decap_8
XFILLER_16_621 VPWR VGND sg13g2_fill_1
XFILLER_44_974 VPWR VGND sg13g2_decap_8
XFILLER_43_462 VPWR VGND sg13g2_fill_1
XFILLER_43_451 VPWR VGND sg13g2_decap_4
XFILLER_15_131 VPWR VGND sg13g2_fill_1
XFILLER_30_145 VPWR VGND sg13g2_fill_1
Xhold308 mydesign.pe_weights\[47\] VPWR VGND net927 sg13g2_dlygate4sd3_1
Xhold319 mydesign.pe_weights\[34\] VPWR VGND net938 sg13g2_dlygate4sd3_1
X_4390_ _1318_ _1308_ _1317_ VPWR VGND sg13g2_xnor2_1
X_3410_ VPWR VGND _0405_ _2698_ _0453_ _0412_ _0456_ _0451_ sg13g2_a221oi_1
X_3341_ net497 _0393_ _0395_ VPWR VGND sg13g2_nor2_2
X_3272_ _2679_ VPWR _0033_ VGND _2520_ _2678_ sg13g2_o21ai_1
X_6060_ net218 VGND VPWR net924 mydesign.accum\[26\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_5011_ _1862_ _1863_ _1864_ VPWR VGND sg13g2_and2_1
XFILLER_19_492 VPWR VGND sg13g2_fill_1
X_5913_ net331 VGND VPWR _0139_ mydesign.pe_weights\[51\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_35_985 VPWR VGND sg13g2_decap_8
X_5844_ net81 VGND VPWR _0070_ net10 clknet_leaf_42_clk sg13g2_dfrbpq_2
XFILLER_22_613 VPWR VGND sg13g2_fill_2
X_5775_ net183 VGND VPWR _0001_ mydesign.weights\[2\]\[4\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_22_679 VPWR VGND sg13g2_decap_8
X_4726_ _1617_ _1618_ _1619_ VPWR VGND sg13g2_nor2b_1
X_4657_ net467 VPWR _1554_ VGND net560 net818 sg13g2_o21ai_1
X_3608_ _0631_ net1004 _0630_ VPWR VGND sg13g2_xnor2_1
X_4588_ _1496_ _1495_ _0209_ VPWR VGND sg13g2_nor2b_1
X_3539_ _0566_ _0565_ _0558_ VPWR VGND sg13g2_nand2b_1
X_5209_ _2039_ _2038_ _2041_ VPWR VGND sg13g2_xor2_1
XFILLER_45_716 VPWR VGND sg13g2_decap_8
XFILLER_26_974 VPWR VGND sg13g2_decap_8
XFILLER_41_944 VPWR VGND sg13g2_decap_8
XFILLER_12_145 VPWR VGND sg13g2_fill_2
XFILLER_16_97 VPWR VGND sg13g2_decap_4
XFILLER_8_138 VPWR VGND sg13g2_fill_2
XFILLER_32_96 VPWR VGND sg13g2_fill_1
XFILLER_48_532 VPWR VGND sg13g2_fill_2
XFILLER_48_565 VPWR VGND sg13g2_fill_2
XFILLER_36_727 VPWR VGND sg13g2_decap_8
XFILLER_36_738 VPWR VGND sg13g2_fill_2
XFILLER_44_771 VPWR VGND sg13g2_decap_8
XFILLER_17_985 VPWR VGND sg13g2_decap_8
XFILLER_31_410 VPWR VGND sg13g2_fill_2
XFILLER_32_922 VPWR VGND sg13g2_decap_8
X_3890_ _0879_ mydesign.accum\[109\] _0878_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_999 VPWR VGND sg13g2_decap_8
X_5560_ _2357_ VPWR _0320_ VGND net603 _2355_ sg13g2_o21ai_1
X_4511_ _1423_ mydesign.pe_weights\[48\] mydesign.pe_inputs\[38\] VPWR VGND sg13g2_nand2_1
X_5491_ _2292_ _2275_ _2294_ VPWR VGND sg13g2_xor2_1
Xhold116 _0272_ VPWR VGND net735 sg13g2_dlygate4sd3_1
Xhold105 _0352_ VPWR VGND net724 sg13g2_dlygate4sd3_1
X_4442_ _1367_ _1365_ _1366_ VPWR VGND sg13g2_nand2_1
Xhold149 mydesign.inputs\[0\]\[21\] VPWR VGND net768 sg13g2_dlygate4sd3_1
Xhold138 mydesign.accum\[108\] VPWR VGND net757 sg13g2_dlygate4sd3_1
Xhold127 _0236_ VPWR VGND net746 sg13g2_dlygate4sd3_1
X_4373_ _1300_ VPWR _1302_ VGND _1298_ _1299_ sg13g2_o21ai_1
X_3324_ _0381_ _0382_ _0059_ VPWR VGND sg13g2_nor2_1
Xfanout618 net619 net618 VPWR VGND sg13g2_buf_8
Xfanout607 net608 net607 VPWR VGND sg13g2_buf_8
Xfanout629 net632 net629 VPWR VGND sg13g2_buf_1
X_6112_ net196 VGND VPWR _0338_ mydesign.out\[2\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_6043_ net286 VGND VPWR net829 mydesign.pe_weights\[17\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3255_ VGND VPWR _2671_ _2657_ _2606_ sg13g2_or2_1
X_3186_ _2622_ _2621_ VPWR VGND sg13g2_inv_2
XFILLER_27_727 VPWR VGND sg13g2_decap_4
XFILLER_23_922 VPWR VGND sg13g2_fill_2
XFILLER_22_421 VPWR VGND sg13g2_fill_2
XFILLER_23_966 VPWR VGND sg13g2_decap_8
X_5827_ net115 VGND VPWR net710 mydesign.inputs\[3\]\[0\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_5758_ net612 VPWR _2509_ VGND net869 _2505_ sg13g2_o21ai_1
X_4709_ _1603_ _1596_ _1601_ VPWR VGND sg13g2_xnor2_1
X_5689_ net457 net456 _2468_ _2470_ VPWR VGND sg13g2_nor3_1
XFILLER_2_804 VPWR VGND sg13g2_decap_8
XFILLER_2_859 VPWR VGND sg13g2_fill_1
XFILLER_18_727 VPWR VGND sg13g2_decap_4
XFILLER_45_546 VPWR VGND sg13g2_fill_2
XFILLER_45_568 VPWR VGND sg13g2_decap_4
XFILLER_41_752 VPWR VGND sg13g2_fill_2
XFILLER_14_977 VPWR VGND sg13g2_decap_8
XFILLER_49_874 VPWR VGND sg13g2_decap_8
X_4991_ _1821_ _1823_ _1843_ _1845_ VPWR VGND sg13g2_or3_1
XFILLER_23_207 VPWR VGND sg13g2_fill_2
XFILLER_23_218 VPWR VGND sg13g2_fill_2
XFILLER_44_590 VPWR VGND sg13g2_fill_1
X_3942_ _0922_ net547 mydesign.weights\[3\]\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_17_1027 VPWR VGND sg13g2_fill_2
X_3873_ _0862_ _0859_ _0863_ VPWR VGND sg13g2_xor2_1
XFILLER_31_262 VPWR VGND sg13g2_decap_4
X_5612_ _2402_ _2387_ _2403_ VPWR VGND sg13g2_xor2_1
XFILLER_20_947 VPWR VGND sg13g2_decap_8
XFILLER_9_970 VPWR VGND sg13g2_decap_8
X_5543_ _2343_ _2325_ _2341_ VPWR VGND sg13g2_xnor2_1
X_5474_ _2277_ net520 mydesign.pe_weights\[20\] VPWR VGND sg13g2_nand2_1
X_5867__39 VPWR VGND net39 sg13g2_tiehi
X_4425_ _1351_ _1345_ _1350_ VPWR VGND sg13g2_nand2_1
X_4356_ net629 VPWR _1291_ VGND mydesign.pe_inputs\[39\] net434 sg13g2_o21ai_1
X_3307_ net742 net429 net618 _2694_ VPWR VGND sg13g2_nand3_1
XFILLER_24_1009 VPWR VGND sg13g2_decap_8
Xfanout437 net438 net437 VPWR VGND sg13g2_buf_8
Xfanout448 net452 net448 VPWR VGND sg13g2_buf_1
X_4287_ VGND VPWR net579 _1228_ _0175_ _1229_ sg13g2_a21oi_1
Xfanout459 _0396_ net459 VPWR VGND sg13g2_buf_8
XFILLER_39_340 VPWR VGND sg13g2_fill_1
X_3238_ _2648_ _2657_ _2658_ VPWR VGND sg13g2_nor2_1
X_6026_ net358 VGND VPWR _0252_ mydesign.pe_inputs\[20\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3169_ _2609_ net1 net432 VPWR VGND sg13g2_nand2_1
X_5832__105 VPWR VGND net105 sg13g2_tiehi
XFILLER_27_513 VPWR VGND sg13g2_fill_1
XFILLER_15_719 VPWR VGND sg13g2_fill_1
XFILLER_27_546 VPWR VGND sg13g2_decap_8
XFILLER_27_557 VPWR VGND sg13g2_fill_1
XFILLER_23_741 VPWR VGND sg13g2_fill_1
XFILLER_22_251 VPWR VGND sg13g2_fill_2
XFILLER_11_947 VPWR VGND sg13g2_decap_8
Xhold480 _0296_ VPWR VGND net1099 sg13g2_dlygate4sd3_1
Xhold491 mydesign.load_counter\[3\] VPWR VGND net1110 sg13g2_dlygate4sd3_1
XFILLER_49_126 VPWR VGND sg13g2_fill_1
XFILLER_18_502 VPWR VGND sg13g2_fill_1
XFILLER_38_62 VPWR VGND sg13g2_decap_4
XFILLER_46_866 VPWR VGND sg13g2_decap_8
XFILLER_45_365 VPWR VGND sg13g2_fill_2
XFILLER_33_527 VPWR VGND sg13g2_fill_1
XFILLER_10_991 VPWR VGND sg13g2_decap_8
Xclkload14 VPWR clkload14/Y clknet_leaf_34_clk VGND sg13g2_inv_1
X_4210_ _1166_ _1164_ _1165_ VPWR VGND sg13g2_xnor2_1
X_5190_ _2023_ net979 _2024_ VPWR VGND sg13g2_xor2_1
X_4141_ _1100_ mydesign.pe_weights\[61\] _1056_ VPWR VGND sg13g2_nand2_1
X_4072_ VGND VPWR net571 _1041_ _0147_ _1042_ sg13g2_a21oi_1
XFILLER_49_671 VPWR VGND sg13g2_decap_8
XFILLER_48_181 VPWR VGND sg13g2_fill_2
XFILLER_24_505 VPWR VGND sg13g2_fill_2
X_4974_ _1829_ _1813_ _1827_ VPWR VGND sg13g2_xnor2_1
X_3925_ _0911_ _2655_ _0910_ VPWR VGND sg13g2_nand2_2
Xclkload8 clkload8/Y clknet_leaf_18_clk VPWR VGND sg13g2_inv_2
X_3856_ _0847_ _0823_ _0846_ VPWR VGND sg13g2_nand2_1
X_3787_ VGND VPWR _2559_ net491 _0120_ _0784_ sg13g2_a21oi_1
X_5526_ _2306_ _2326_ _2327_ VPWR VGND sg13g2_nor2b_1
X_5457_ _2261_ mydesign.pe_inputs\[9\] mydesign.pe_weights\[21\] VPWR VGND sg13g2_nand2_1
X_4408_ _1333_ _1326_ _1335_ VPWR VGND sg13g2_xor2_1
X_5388_ _2202_ _2200_ _2201_ VPWR VGND sg13g2_nand2_1
X_4339_ _1277_ VPWR _1279_ VGND _1261_ _1264_ sg13g2_o21ai_1
X_5953__251 VPWR VGND net251 sg13g2_tiehi
XFILLER_46_118 VPWR VGND sg13g2_fill_2
XFILLER_46_107 VPWR VGND sg13g2_fill_1
X_6009_ net54 VGND VPWR net790 mydesign.pe_weights\[27\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_43_858 VPWR VGND sg13g2_decap_8
XFILLER_15_549 VPWR VGND sg13g2_decap_4
XFILLER_11_700 VPWR VGND sg13g2_fill_2
XFILLER_23_560 VPWR VGND sg13g2_fill_1
X_6129__372 VPWR VGND net372 sg13g2_tiehi
XFILLER_23_582 VPWR VGND sg13g2_decap_4
XFILLER_40_63 VPWR VGND sg13g2_decap_8
XFILLER_46_1020 VPWR VGND sg13g2_decap_8
XFILLER_49_50 VPWR VGND sg13g2_decap_4
X_6032__330 VPWR VGND net330 sg13g2_tiehi
XFILLER_46_663 VPWR VGND sg13g2_decap_8
XFILLER_34_825 VPWR VGND sg13g2_fill_1
XFILLER_33_379 VPWR VGND sg13g2_decap_8
XFILLER_42_891 VPWR VGND sg13g2_decap_8
XFILLER_14_560 VPWR VGND sg13g2_fill_2
X_3710_ _0719_ _0711_ _0720_ VPWR VGND sg13g2_xor2_1
XFILLER_14_1019 VPWR VGND sg13g2_decap_8
X_4690_ _1585_ _1560_ _1584_ VPWR VGND sg13g2_nand2_1
X_3641_ _0656_ net545 net555 mydesign.weights\[1\]\[15\] VPWR VGND sg13g2_and3_1
X_3572_ _0596_ _0597_ _0092_ VPWR VGND sg13g2_nor2_1
X_5311_ _2134_ VPWR _0294_ VGND net599 _2130_ sg13g2_o21ai_1
X_5242_ _2073_ _2051_ _2072_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
X_5173_ VPWR _2010_ _2009_ VGND sg13g2_inv_1
X_4124_ _1081_ _1082_ _1083_ _1084_ VPWR VGND sg13g2_nor3_1
XFILLER_29_619 VPWR VGND sg13g2_fill_2
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_2
X_4055_ _1010_ VPWR _1027_ VGND _1009_ _1012_ sg13g2_o21ai_1
Xclkbuf_leaf_48_clk clknet_3_1__leaf_clk clknet_leaf_48_clk VPWR VGND sg13g2_buf_8
XFILLER_12_519 VPWR VGND sg13g2_decap_8
XFILLER_24_346 VPWR VGND sg13g2_fill_1
X_4957_ _1808_ VPWR _1812_ VGND _1794_ _1809_ sg13g2_o21ai_1
X_4888_ net623 _1761_ _1762_ VPWR VGND sg13g2_and2_1
X_3908_ VGND VPWR mydesign.accum\[109\] _0878_ _0896_ _0880_ sg13g2_a21oi_1
X_3839_ VGND VPWR _0831_ _0830_ _0815_ sg13g2_or2_1
X_5509_ _2309_ _2308_ _2311_ VPWR VGND sg13g2_xor2_1
XFILLER_0_957 VPWR VGND sg13g2_decap_8
X_5836__97 VPWR VGND net97 sg13g2_tiehi
Xclkbuf_leaf_39_clk clknet_3_4__leaf_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_43_644 VPWR VGND sg13g2_fill_2
XFILLER_43_633 VPWR VGND sg13g2_decap_8
XFILLER_37_1008 VPWR VGND sg13g2_decap_8
XFILLER_11_574 VPWR VGND sg13g2_decap_4
XFILLER_7_578 VPWR VGND sg13g2_fill_1
XFILLER_39_928 VPWR VGND sg13g2_decap_8
XFILLER_38_405 VPWR VGND sg13g2_decap_8
XFILLER_47_950 VPWR VGND sg13g2_decap_8
XFILLER_38_449 VPWR VGND sg13g2_decap_8
X_5860_ net53 VGND VPWR _0086_ mydesign.pe_weights\[62\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_4811_ _1690_ _1688_ _1689_ VPWR VGND sg13g2_nand2_1
X_5791_ net159 VGND VPWR _0017_ mydesign.inputs\[2\]\[4\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_6108__220 VPWR VGND net220 sg13g2_tiehi
X_4742_ _1614_ _1618_ _1634_ VPWR VGND sg13g2_and2_1
X_4673_ _1569_ _1552_ _1567_ VPWR VGND sg13g2_xnor2_1
X_3624_ VGND VPWR _0640_ _0641_ _0642_ net542 sg13g2_a21oi_1
X_3555_ _0581_ _0506_ _0523_ VPWR VGND sg13g2_nand2_1
X_3486_ net553 mydesign.weights\[0\]\[25\] mydesign.weights\[0\]\[21\] mydesign.weights\[0\]\[17\]
+ mydesign.weights\[0\]\[13\] net546 _0519_ VPWR VGND sg13g2_mux4_1
X_5225_ _2009_ mydesign.pe_weights\[30\] _2056_ VPWR VGND sg13g2_nor2b_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
X_5156_ _1995_ net889 _1981_ VPWR VGND sg13g2_xnor2_1
X_4107_ _1068_ net1003 _1069_ VPWR VGND sg13g2_xor2_1
X_5087_ _1908_ _1929_ _1930_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_972 VPWR VGND sg13g2_decap_8
X_4038_ net428 mydesign.pe_inputs\[54\] mydesign.accum\[101\] _1011_ VPWR VGND sg13g2_a21o_1
XFILLER_37_482 VPWR VGND sg13g2_fill_1
XFILLER_40_614 VPWR VGND sg13g2_fill_2
X_5989_ net170 VGND VPWR _0215_ mydesign.pe_inputs\[31\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_4_515 VPWR VGND sg13g2_fill_2
X_5805__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_0_732 VPWR VGND sg13g2_decap_8
XFILLER_43_1012 VPWR VGND sg13g2_decap_8
XFILLER_0_743 VPWR VGND sg13g2_fill_2
XFILLER_48_769 VPWR VGND sg13g2_decap_8
XFILLER_47_235 VPWR VGND sg13g2_fill_2
XFILLER_36_909 VPWR VGND sg13g2_decap_8
XFILLER_29_972 VPWR VGND sg13g2_decap_8
XFILLER_28_482 VPWR VGND sg13g2_decap_8
XFILLER_44_953 VPWR VGND sg13g2_decap_8
XFILLER_31_614 VPWR VGND sg13g2_fill_2
XFILLER_12_861 VPWR VGND sg13g2_fill_1
XFILLER_8_865 VPWR VGND sg13g2_decap_4
XFILLER_12_894 VPWR VGND sg13g2_fill_2
XFILLER_7_375 VPWR VGND sg13g2_decap_4
Xhold309 mydesign.accum\[9\] VPWR VGND net928 sg13g2_dlygate4sd3_1
X_3340_ net544 net554 _0394_ VPWR VGND sg13g2_and2_1
X_3271_ net617 _2678_ net670 _2679_ VPWR VGND sg13g2_nand3_1
X_5010_ _1840_ _1842_ _1861_ _1863_ VPWR VGND sg13g2_or3_1
XFILLER_39_758 VPWR VGND sg13g2_decap_8
XFILLER_26_408 VPWR VGND sg13g2_fill_2
X_5912_ net333 VGND VPWR _0138_ mydesign.pe_weights\[50\] clknet_leaf_45_clk sg13g2_dfrbpq_2
XFILLER_35_964 VPWR VGND sg13g2_decap_8
X_5843_ net83 VGND VPWR net1070 net9 clknet_leaf_43_clk sg13g2_dfrbpq_2
XFILLER_22_603 VPWR VGND sg13g2_fill_2
X_5774_ net240 VGND VPWR _0000_ mydesign.valid_out clknet_leaf_49_clk sg13g2_dfrbpq_1
XFILLER_21_168 VPWR VGND sg13g2_fill_2
X_4725_ _1537_ _1616_ mydesign.pe_weights\[46\] _1618_ VPWR VGND sg13g2_nand3_1
X_4656_ _1551_ _1550_ _1553_ VPWR VGND sg13g2_xor2_1
X_3607_ _0616_ VPWR _0630_ VGND _0615_ _0617_ sg13g2_o21ai_1
X_4587_ net473 VPWR _1496_ VGND net574 net861 sg13g2_o21ai_1
X_3538_ _0565_ _0541_ _0563_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_1018 VPWR VGND sg13g2_decap_8
X_3469_ _0505_ _0394_ mydesign.inputs\[0\]\[14\] net495 mydesign.inputs\[0\]\[18\]
+ VPWR VGND sg13g2_a22oi_1
X_5208_ _2038_ _2039_ _2040_ VPWR VGND sg13g2_nor2_1
X_5139_ net475 VPWR _1980_ VGND net584 net1005 sg13g2_o21ai_1
XFILLER_29_213 VPWR VGND sg13g2_decap_8
XFILLER_44_216 VPWR VGND sg13g2_fill_1
XFILLER_26_953 VPWR VGND sg13g2_decap_8
XFILLER_41_923 VPWR VGND sg13g2_decap_8
XFILLER_16_54 VPWR VGND sg13g2_fill_1
XFILLER_25_474 VPWR VGND sg13g2_fill_1
XFILLER_40_433 VPWR VGND sg13g2_fill_2
XFILLER_40_477 VPWR VGND sg13g2_decap_8
XFILLER_8_106 VPWR VGND sg13g2_decap_4
XFILLER_21_680 VPWR VGND sg13g2_fill_1
XFILLER_32_86 VPWR VGND sg13g2_fill_1
XFILLER_5_835 VPWR VGND sg13g2_fill_1
XFILLER_4_334 VPWR VGND sg13g2_fill_1
XFILLER_4_378 VPWR VGND sg13g2_fill_2
XFILLER_35_227 VPWR VGND sg13g2_fill_2
XFILLER_44_750 VPWR VGND sg13g2_decap_8
XFILLER_17_964 VPWR VGND sg13g2_decap_8
XFILLER_32_901 VPWR VGND sg13g2_decap_8
XFILLER_43_271 VPWR VGND sg13g2_fill_2
X_6029__346 VPWR VGND net346 sg13g2_tiehi
XFILLER_31_477 VPWR VGND sg13g2_fill_1
XFILLER_32_978 VPWR VGND sg13g2_decap_8
XFILLER_31_499 VPWR VGND sg13g2_fill_2
XFILLER_8_673 VPWR VGND sg13g2_decap_8
X_4510_ VGND VPWR net574 _1421_ _0205_ _1422_ sg13g2_a21oi_1
X_5490_ _2292_ _2275_ _2293_ VPWR VGND sg13g2_nor2b_1
Xhold106 mydesign.weights\[3\]\[0\] VPWR VGND net725 sg13g2_dlygate4sd3_1
Xhold117 mydesign.inputs\[2\]\[19\] VPWR VGND net736 sg13g2_dlygate4sd3_1
X_4441_ mydesign.pe_inputs\[42\] mydesign.pe_weights\[55\] mydesign.accum\[77\] _1366_
+ VPWR VGND sg13g2_a21o_1
Xhold128 mydesign.weights\[2\]\[4\] VPWR VGND net747 sg13g2_dlygate4sd3_1
Xhold139 mydesign.accum\[16\] VPWR VGND net758 sg13g2_dlygate4sd3_1
X_4372_ _1298_ _1299_ _1300_ _1301_ VPWR VGND sg13g2_nor3_1
X_6111_ net204 VGND VPWR _0337_ mydesign.out\[1\] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_3323_ _0382_ net614 _0380_ VPWR VGND sg13g2_nand2_1
Xfanout608 net609 net608 VPWR VGND sg13g2_buf_8
Xfanout619 net640 net619 VPWR VGND sg13g2_buf_8
X_3254_ net800 _2670_ _2659_ _0024_ VPWR VGND sg13g2_mux2_1
X_6042_ net290 VGND VPWR net904 mydesign.pe_weights\[16\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3185_ mydesign.load_counter\[3\] net596 _2621_ VPWR VGND sg13g2_nor2_1
X_5912__333 VPWR VGND net333 sg13g2_tiehi
X_5826_ net116 VGND VPWR _0052_ mydesign.inputs\[0\]\[19\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5757_ VGND VPWR _1773_ _2505_ _0366_ net931 sg13g2_a21oi_1
XFILLER_10_639 VPWR VGND sg13g2_decap_8
XFILLER_33_1022 VPWR VGND sg13g2_decap_8
X_4708_ _1596_ _1601_ _1602_ VPWR VGND sg13g2_and2_1
X_5688_ _2469_ VPWR _0336_ VGND net755 _2468_ sg13g2_o21ai_1
X_4639_ net624 VPWR _1540_ VGND mydesign.pe_weights\[29\] net437 sg13g2_o21ai_1
XFILLER_2_849 VPWR VGND sg13g2_fill_2
XFILLER_1_359 VPWR VGND sg13g2_decap_4
XFILLER_40_1015 VPWR VGND sg13g2_decap_8
XFILLER_27_86 VPWR VGND sg13g2_decap_8
XFILLER_14_912 VPWR VGND sg13g2_fill_2
XFILLER_41_720 VPWR VGND sg13g2_decap_8
X_5887__376 VPWR VGND net376 sg13g2_tiehi
XFILLER_14_956 VPWR VGND sg13g2_decap_8
X_5963__231 VPWR VGND net231 sg13g2_tiehi
XFILLER_5_621 VPWR VGND sg13g2_decap_4
XFILLER_0_370 VPWR VGND sg13g2_fill_1
XFILLER_49_853 VPWR VGND sg13g2_decap_8
XFILLER_1_1020 VPWR VGND sg13g2_decap_8
X_4990_ _1843_ VPWR _1844_ VGND _1821_ _1823_ sg13g2_o21ai_1
X_3941_ _0921_ mydesign.weights\[3\]\[10\] net547 VPWR VGND sg13g2_nand2b_1
XFILLER_17_1006 VPWR VGND sg13g2_decap_8
XFILLER_32_720 VPWR VGND sg13g2_fill_2
X_3872_ _0862_ _0860_ _0861_ VPWR VGND sg13g2_nand2_1
XFILLER_20_926 VPWR VGND sg13g2_decap_8
X_5611_ _2402_ _2388_ _2400_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_797 VPWR VGND sg13g2_decap_4
X_5542_ _2324_ _2341_ _2323_ _2342_ VPWR VGND sg13g2_nand3_1
XFILLER_8_481 VPWR VGND sg13g2_fill_1
X_5473_ _2267_ VPWR _2276_ VGND _2260_ _2268_ sg13g2_o21ai_1
X_4424_ _1349_ _1346_ _1350_ VPWR VGND sg13g2_xor2_1
X_4355_ VGND VPWR _2561_ net434 _0182_ _1290_ sg13g2_a21oi_1
X_3306_ _2693_ VPWR _0053_ VGND net603 net429 sg13g2_o21ai_1
Xfanout438 net439 net438 VPWR VGND sg13g2_buf_8
X_4286_ net471 VPWR _1229_ VGND net579 net911 sg13g2_o21ai_1
Xfanout449 net450 net449 VPWR VGND sg13g2_buf_8
X_6025_ net362 VGND VPWR net822 mydesign.weights\[3\]\[11\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3237_ _2657_ _2588_ net596 VPWR VGND sg13g2_nand2_2
X_3168_ _2605_ _2606_ _2607_ _2608_ VPWR VGND sg13g2_nor3_1
XFILLER_27_536 VPWR VGND sg13g2_fill_2
XFILLER_39_396 VPWR VGND sg13g2_decap_8
X_3099_ VPWR _2540_ net528 VGND sg13g2_inv_1
XFILLER_42_539 VPWR VGND sg13g2_decap_8
XFILLER_23_775 VPWR VGND sg13g2_fill_1
X_5809_ net135 VGND VPWR _0035_ mydesign.inputs\[2\]\[18\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_13_55 VPWR VGND sg13g2_fill_1
XFILLER_22_296 VPWR VGND sg13g2_decap_8
Xhold481 mydesign.pe_inputs\[44\] VPWR VGND net1100 sg13g2_dlygate4sd3_1
Xhold470 mydesign.accum\[13\] VPWR VGND net1089 sg13g2_dlygate4sd3_1
Xhold492 mydesign.pe_inputs\[4\] VPWR VGND net1111 sg13g2_dlygate4sd3_1
XFILLER_38_41 VPWR VGND sg13g2_fill_1
XFILLER_45_311 VPWR VGND sg13g2_fill_2
XFILLER_46_845 VPWR VGND sg13g2_decap_8
XFILLER_18_536 VPWR VGND sg13g2_decap_8
XFILLER_41_550 VPWR VGND sg13g2_fill_1
XFILLER_13_241 VPWR VGND sg13g2_fill_2
XFILLER_9_234 VPWR VGND sg13g2_fill_1
Xclkload15 VPWR clkload15/Y clknet_leaf_37_clk VGND sg13g2_inv_1
XFILLER_10_970 VPWR VGND sg13g2_decap_8
X_5783__171 VPWR VGND net171 sg13g2_tiehi
X_5998__102 VPWR VGND net102 sg13g2_tiehi
X_4140_ VPWR _1099_ _1098_ VGND sg13g2_inv_1
XFILLER_49_650 VPWR VGND sg13g2_decap_8
X_4071_ net464 VPWR _1042_ VGND net566 net940 sg13g2_o21ai_1
XFILLER_37_823 VPWR VGND sg13g2_fill_2
XFILLER_37_889 VPWR VGND sg13g2_decap_8
X_4973_ _1813_ _1827_ _1828_ VPWR VGND sg13g2_and2_1
X_3924_ net615 VPWR _0910_ VGND _2622_ _2683_ sg13g2_o21ai_1
X_6146__164 VPWR VGND net164 sg13g2_tiehi
XFILLER_20_734 VPWR VGND sg13g2_fill_2
Xclkload9 clkload9/Y clknet_leaf_20_clk VPWR VGND sg13g2_inv_2
X_3855_ _0846_ _0837_ _0844_ VPWR VGND sg13g2_xnor2_1
X_3786_ net629 VPWR _0784_ VGND net491 _0783_ sg13g2_o21ai_1
XFILLER_20_789 VPWR VGND sg13g2_fill_1
XFILLER_30_1025 VPWR VGND sg13g2_decap_4
X_5525_ _2324_ _2323_ _2326_ VPWR VGND sg13g2_xor2_1
X_5456_ _2260_ mydesign.pe_inputs\[10\] mydesign.pe_weights\[20\] VPWR VGND sg13g2_nand2_1
X_4407_ _1326_ _1333_ _1334_ VPWR VGND sg13g2_nor2_1
XFILLER_8_1015 VPWR VGND sg13g2_decap_8
X_5387_ _2180_ VPWR _2201_ VGND _2169_ _2181_ sg13g2_o21ai_1
X_4338_ _1261_ _1264_ _1277_ _1278_ VPWR VGND sg13g2_nor3_1
X_5848__73 VPWR VGND net73 sg13g2_tiehi
X_4269_ _1212_ mydesign.pe_weights\[57\] mydesign.pe_inputs\[46\] VPWR VGND sg13g2_nand2_1
X_6008_ net58 VGND VPWR net814 mydesign.pe_weights\[26\] clknet_leaf_26_clk sg13g2_dfrbpq_2
XFILLER_28_867 VPWR VGND sg13g2_decap_8
XFILLER_43_837 VPWR VGND sg13g2_decap_8
XFILLER_42_325 VPWR VGND sg13g2_fill_1
XFILLER_11_789 VPWR VGND sg13g2_fill_1
XFILLER_40_97 VPWR VGND sg13g2_fill_1
XFILLER_3_999 VPWR VGND sg13g2_decap_8
XFILLER_2_498 VPWR VGND sg13g2_fill_2
X_5854__65 VPWR VGND net65 sg13g2_tiehi
XFILLER_46_642 VPWR VGND sg13g2_decap_8
XFILLER_18_355 VPWR VGND sg13g2_fill_2
XFILLER_33_314 VPWR VGND sg13g2_decap_8
XFILLER_42_870 VPWR VGND sg13g2_decap_8
XFILLER_14_583 VPWR VGND sg13g2_fill_2
X_3640_ mydesign.weights\[1\]\[11\] net460 net498 _0655_ VPWR VGND sg13g2_nand3_1
X_3571_ net468 VPWR _0597_ VGND net559 net1079 sg13g2_o21ai_1
X_5310_ _2134_ net427 _2131_ VPWR VGND sg13g2_nand2_1
XFILLER_5_292 VPWR VGND sg13g2_fill_1
X_5241_ _2072_ _2052_ _2069_ VPWR VGND sg13g2_xnor2_1
X_5172_ VPWR VGND mydesign.inputs\[3\]\[13\] _2008_ _0395_ mydesign.inputs\[3\]\[1\]
+ _2009_ net454 sg13g2_a221oi_1
X_4123_ _1083_ mydesign.pe_weights\[61\] _1051_ VPWR VGND sg13g2_nand2_1
X_4054_ _1026_ _1025_ _1024_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_119 VPWR VGND sg13g2_decap_8
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_2
XFILLER_37_653 VPWR VGND sg13g2_fill_1
XFILLER_24_314 VPWR VGND sg13g2_decap_8
XFILLER_25_848 VPWR VGND sg13g2_fill_2
X_6007__62 VPWR VGND net62 sg13g2_tiehi
X_4956_ VGND VPWR net589 _1810_ _0262_ _1811_ sg13g2_a21oi_1
X_5909__338 VPWR VGND net338 sg13g2_tiehi
X_4887_ _2606_ _2607_ _2618_ _1761_ VPWR VGND sg13g2_or3_1
XFILLER_20_520 VPWR VGND sg13g2_fill_1
XFILLER_20_542 VPWR VGND sg13g2_fill_2
X_3907_ _0895_ _0894_ _0893_ VPWR VGND sg13g2_nand2b_1
X_3838_ _0830_ _0812_ _0828_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_719 VPWR VGND sg13g2_fill_2
X_3769_ _0773_ net701 _0770_ VPWR VGND sg13g2_nand2_1
X_5508_ _2310_ _2308_ _2309_ VPWR VGND sg13g2_nand2_1
X_5439_ VGND VPWR _2522_ net444 _0310_ _2246_ sg13g2_a21oi_1
XFILLER_0_936 VPWR VGND sg13g2_decap_8
XFILLER_28_631 VPWR VGND sg13g2_decap_8
X_5851__68 VPWR VGND net68 sg13g2_tiehi
XFILLER_16_859 VPWR VGND sg13g2_fill_1
X_5988__178 VPWR VGND net178 sg13g2_tiehi
XFILLER_42_188 VPWR VGND sg13g2_fill_2
XFILLER_24_870 VPWR VGND sg13g2_fill_1
XFILLER_7_557 VPWR VGND sg13g2_decap_4
X_5780__174 VPWR VGND net174 sg13g2_tiehi
XFILLER_2_251 VPWR VGND sg13g2_decap_4
XFILLER_39_907 VPWR VGND sg13g2_decap_8
XFILLER_38_428 VPWR VGND sg13g2_fill_1
XFILLER_20_1024 VPWR VGND sg13g2_decap_4
XFILLER_46_494 VPWR VGND sg13g2_decap_8
X_4810_ mydesign.pe_inputs\[28\] net533 mydesign.accum\[51\] _1689_ VPWR VGND sg13g2_a21o_1
X_5790_ net160 VGND VPWR net643 mydesign.inputs\[2\]\[11\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_4741_ _1633_ _1632_ _1631_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_862 VPWR VGND sg13g2_fill_2
X_4672_ VGND VPWR _1568_ _1567_ _1552_ sg13g2_or2_1
X_3623_ _0641_ _0394_ mydesign.weights\[1\]\[12\] net461 mydesign.weights\[1\]\[20\]
+ VPWR VGND sg13g2_a22oi_1
X_3554_ _0561_ VPWR _0580_ VGND _0559_ _0562_ sg13g2_o21ai_1
X_3485_ VGND VPWR _2578_ net484 _0084_ _0518_ sg13g2_a21oi_1
X_5224_ mydesign.pe_weights\[29\] _2015_ _2055_ VPWR VGND sg13g2_and2_1
XFILLER_5_1007 VPWR VGND sg13g2_decap_8
X_5155_ VGND VPWR _1970_ _1985_ _1994_ _1984_ sg13g2_a21oi_1
X_4106_ _1068_ net561 _1067_ VPWR VGND sg13g2_nand2_1
XFILLER_38_951 VPWR VGND sg13g2_decap_8
X_5086_ _1928_ _1925_ _1929_ VPWR VGND sg13g2_xor2_1
XFILLER_37_461 VPWR VGND sg13g2_decap_8
XFILLER_37_450 VPWR VGND sg13g2_fill_2
X_4037_ mydesign.pe_inputs\[54\] net428 mydesign.accum\[101\] _1010_ VPWR VGND sg13g2_nand3_1
XFILLER_37_472 VPWR VGND sg13g2_fill_2
XFILLER_13_818 VPWR VGND sg13g2_fill_1
XFILLER_24_177 VPWR VGND sg13g2_fill_2
X_5988_ net178 VGND VPWR _0214_ mydesign.pe_inputs\[30\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_4939_ net477 VPWR _1796_ VGND net585 net949 sg13g2_o21ai_1
XFILLER_21_851 VPWR VGND sg13g2_fill_1
X_5922__313 VPWR VGND net313 sg13g2_tiehi
XFILLER_21_895 VPWR VGND sg13g2_decap_8
X_6133__336 VPWR VGND net336 sg13g2_tiehi
XFILLER_48_748 VPWR VGND sg13g2_decap_8
XFILLER_29_951 VPWR VGND sg13g2_decap_8
XFILLER_35_409 VPWR VGND sg13g2_decap_8
XFILLER_44_932 VPWR VGND sg13g2_decap_8
XFILLER_15_100 VPWR VGND sg13g2_decap_8
XFILLER_43_442 VPWR VGND sg13g2_decap_4
XFILLER_43_420 VPWR VGND sg13g2_decap_4
XFILLER_15_166 VPWR VGND sg13g2_fill_2
XFILLER_31_659 VPWR VGND sg13g2_fill_1
X_3270_ _2678_ _2663_ VPWR VGND _2662_ sg13g2_nand2b_2
X_5973__211 VPWR VGND net211 sg13g2_tiehi
XFILLER_30_5 VPWR VGND sg13g2_fill_2
X_5911_ net335 VGND VPWR _0137_ mydesign.pe_weights\[49\] clknet_leaf_45_clk sg13g2_dfrbpq_2
XFILLER_35_943 VPWR VGND sg13g2_decap_8
X_5842_ net85 VGND VPWR _0068_ net8 clknet_leaf_7_clk sg13g2_dfrbpq_2
XFILLER_22_659 VPWR VGND sg13g2_decap_8
X_5773_ _2515_ VPWR _0375_ VGND net598 _2511_ sg13g2_o21ai_1
X_4724_ VGND VPWR mydesign.pe_weights\[46\] _1537_ _1617_ _1616_ sg13g2_a21oi_1
XFILLER_30_670 VPWR VGND sg13g2_decap_8
X_4655_ net815 _1521_ net686 _1552_ VPWR VGND _1550_ sg13g2_nand4_1
X_3606_ _0629_ _0623_ _0626_ VPWR VGND sg13g2_nand2_1
X_4586_ net574 VPWR _1495_ VGND _1493_ _1494_ sg13g2_o21ai_1
X_3537_ _0564_ _0563_ _0541_ VPWR VGND sg13g2_nand2b_1
X_3468_ VGND VPWR net554 mydesign.inputs\[0\]\[22\] _0504_ _0503_ sg13g2_a21oi_1
X_3399_ VGND VPWR _0445_ _0446_ net517 mydesign.accum\[3\] sg13g2_a21oi_2
X_5207_ _2039_ mydesign.pe_weights\[29\] _2010_ VPWR VGND sg13g2_nand2_1
XFILLER_29_203 VPWR VGND sg13g2_decap_4
X_5138_ net584 VPWR _1979_ VGND _1977_ _1978_ sg13g2_o21ai_1
XFILLER_17_409 VPWR VGND sg13g2_fill_2
XFILLER_38_781 VPWR VGND sg13g2_fill_2
X_5069_ _1913_ _1896_ _1912_ VPWR VGND sg13g2_nand2_1
XFILLER_41_902 VPWR VGND sg13g2_decap_8
XFILLER_41_979 VPWR VGND sg13g2_decap_8
XFILLER_12_158 VPWR VGND sg13g2_fill_1
XFILLER_4_313 VPWR VGND sg13g2_fill_2
XFILLER_10_1012 VPWR VGND sg13g2_decap_8
XFILLER_0_552 VPWR VGND sg13g2_fill_2
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_48_567 VPWR VGND sg13g2_fill_1
XFILLER_17_943 VPWR VGND sg13g2_decap_8
XFILLER_28_291 VPWR VGND sg13g2_decap_8
XFILLER_43_294 VPWR VGND sg13g2_decap_8
XFILLER_16_497 VPWR VGND sg13g2_fill_1
XFILLER_31_412 VPWR VGND sg13g2_fill_1
XFILLER_32_957 VPWR VGND sg13g2_decap_8
XFILLER_31_456 VPWR VGND sg13g2_fill_2
XFILLER_12_681 VPWR VGND sg13g2_decap_4
XFILLER_11_180 VPWR VGND sg13g2_fill_2
Xhold107 _0340_ VPWR VGND net726 sg13g2_dlygate4sd3_1
X_4440_ mydesign.pe_weights\[55\] mydesign.pe_inputs\[42\] mydesign.accum\[77\] _1365_
+ VPWR VGND sg13g2_nand3_1
Xhold129 mydesign.weights\[0\]\[16\] VPWR VGND net748 sg13g2_dlygate4sd3_1
Xhold118 mydesign.weights\[1\]\[22\] VPWR VGND net737 sg13g2_dlygate4sd3_1
XFILLER_4_880 VPWR VGND sg13g2_decap_4
X_4371_ _1300_ mydesign.pe_weights\[52\] mydesign.pe_inputs\[41\] VPWR VGND sg13g2_nand2_1
X_6110_ net212 VGND VPWR _0336_ mydesign.out\[0\] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_3322_ VGND VPWR _2600_ _2647_ _0381_ net596 sg13g2_a21oi_1
Xfanout609 _2590_ net609 VPWR VGND sg13g2_buf_8
X_3253_ net4 _2666_ _2670_ VPWR VGND sg13g2_and2_1
X_6041_ net294 VGND VPWR _0267_ mydesign.accum\[47\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_3184_ VPWR _2620_ _2619_ VGND sg13g2_inv_1
XFILLER_14_0 VPWR VGND sg13g2_fill_2
X_5825_ net117 VGND VPWR _0051_ mydesign.inputs\[0\]\[18\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_33_1001 VPWR VGND sg13g2_decap_8
X_5756_ net612 VPWR _2508_ VGND net930 _2505_ sg13g2_o21ai_1
X_5687_ _2469_ net755 _2466_ VPWR VGND sg13g2_nand2_1
X_4707_ _1600_ _1597_ _1601_ VPWR VGND sg13g2_xor2_1
X_4638_ VGND VPWR _2552_ net439 _0216_ _1539_ sg13g2_a21oi_1
X_4569_ _1477_ _1478_ _0208_ VPWR VGND sg13g2_nor2_1
XFILLER_1_316 VPWR VGND sg13g2_decap_4
XFILLER_45_526 VPWR VGND sg13g2_fill_2
XFILLER_45_515 VPWR VGND sg13g2_fill_2
XFILLER_32_209 VPWR VGND sg13g2_fill_1
XFILLER_40_220 VPWR VGND sg13g2_decap_4
XFILLER_14_935 VPWR VGND sg13g2_decap_8
XFILLER_25_261 VPWR VGND sg13g2_decap_4
XFILLER_26_795 VPWR VGND sg13g2_decap_8
XFILLER_41_754 VPWR VGND sg13g2_fill_1
XFILLER_13_445 VPWR VGND sg13g2_fill_2
XFILLER_40_275 VPWR VGND sg13g2_fill_1
XFILLER_5_655 VPWR VGND sg13g2_decap_4
XFILLER_1_861 VPWR VGND sg13g2_fill_1
XFILLER_49_832 VPWR VGND sg13g2_decap_8
XFILLER_1_894 VPWR VGND sg13g2_decap_8
X_5777__179 VPWR VGND net179 sg13g2_tiehi
XFILLER_48_353 VPWR VGND sg13g2_fill_2
XFILLER_36_559 VPWR VGND sg13g2_fill_2
X_3940_ VGND VPWR _2555_ net486 _0137_ _0920_ sg13g2_a21oi_1
X_3871_ _0804_ mydesign.pe_inputs\[57\] mydesign.accum\[108\] _0861_ VPWR VGND sg13g2_a21o_1
X_5610_ _2401_ _2388_ _2400_ VPWR VGND sg13g2_nand2_1
XFILLER_31_275 VPWR VGND sg13g2_fill_2
X_5541_ _2339_ _2340_ _2341_ VPWR VGND sg13g2_and2_1
XFILLER_8_460 VPWR VGND sg13g2_decap_8
X_5472_ _2271_ VPWR _2275_ VGND _2257_ _2272_ sg13g2_o21ai_1
X_4423_ _1349_ _1347_ _1348_ VPWR VGND sg13g2_nand2_1
X_4354_ net628 VPWR _1290_ VGND mydesign.pe_inputs\[38\] net434 sg13g2_o21ai_1
Xfanout428 _0933_ net428 VPWR VGND sg13g2_buf_8
X_3305_ net709 net429 net618 _2693_ VPWR VGND sg13g2_nand3_1
Xfanout439 net453 net439 VPWR VGND sg13g2_buf_8
X_4285_ _1226_ _1209_ _1228_ VPWR VGND sg13g2_xor2_1
X_6024_ net366 VGND VPWR net855 mydesign.weights\[3\]\[10\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3236_ net596 _2647_ _2656_ VPWR VGND sg13g2_and2_1
X_3167_ _2607_ mydesign.load_counter\[3\] net596 VPWR VGND sg13g2_nand2_2
XFILLER_27_526 VPWR VGND sg13g2_decap_4
X_3098_ VPWR _2539_ net849 VGND sg13g2_inv_1
XFILLER_42_518 VPWR VGND sg13g2_fill_1
X_5808_ net137 VGND VPWR _0034_ mydesign.inputs\[2\]\[17\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_6_408 VPWR VGND sg13g2_fill_1
X_5739_ _2498_ VPWR _0358_ VGND net600 _2495_ sg13g2_o21ai_1
Xhold460 mydesign.accum\[124\] VPWR VGND net1079 sg13g2_dlygate4sd3_1
Xhold471 mydesign.pe_inputs\[30\] VPWR VGND net1090 sg13g2_dlygate4sd3_1
X_5866__41 VPWR VGND net41 sg13g2_tiehi
Xhold482 mydesign.pe_weights\[39\] VPWR VGND net1101 sg13g2_dlygate4sd3_1
X_6122__56 VPWR VGND net56 sg13g2_tiehi
XFILLER_46_824 VPWR VGND sg13g2_decap_8
XFILLER_45_367 VPWR VGND sg13g2_fill_1
X_5930__297 VPWR VGND net297 sg13g2_tiehi
Xclkload16 clkload16/Y clknet_leaf_31_clk VPWR VGND sg13g2_inv_2
XFILLER_6_986 VPWR VGND sg13g2_decap_8
X_4070_ _1041_ _1037_ _1040_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_1022 VPWR VGND sg13g2_decap_8
XFILLER_17_581 VPWR VGND sg13g2_fill_1
X_4972_ _1826_ _1814_ _1827_ VPWR VGND sg13g2_xor2_1
XFILLER_36_389 VPWR VGND sg13g2_decap_8
X_3923_ VGND VPWR net578 _0908_ _0131_ _0909_ sg13g2_a21oi_1
X_3854_ _0845_ _0844_ _0837_ VPWR VGND sg13g2_nand2b_1
X_5981__195 VPWR VGND net195 sg13g2_tiehi
X_3785_ _0780_ VPWR _0783_ VGND _0781_ _0782_ sg13g2_o21ai_1
XFILLER_30_1004 VPWR VGND sg13g2_decap_8
XFILLER_8_290 VPWR VGND sg13g2_fill_1
X_5524_ _2325_ _2323_ _2324_ VPWR VGND sg13g2_nand2_1
X_5455_ VGND VPWR net588 _2258_ _0313_ _2259_ sg13g2_a21oi_1
X_4406_ _1331_ _1310_ _1333_ VPWR VGND sg13g2_xor2_1
X_5386_ _2198_ _2199_ _2200_ VPWR VGND sg13g2_and2_1
X_4337_ _1277_ _1259_ _1275_ VPWR VGND sg13g2_xnor2_1
X_4268_ _1211_ mydesign.pe_weights\[56\] mydesign.pe_inputs\[47\] VPWR VGND sg13g2_nand2_1
XFILLER_39_150 VPWR VGND sg13g2_fill_1
X_3219_ _2645_ net667 _2642_ VPWR VGND sg13g2_nand2_1
X_6007_ net62 VGND VPWR net857 mydesign.pe_weights\[25\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_4199_ VPWR VGND _1155_ net462 _1154_ net500 _0161_ _2573_ sg13g2_a221oi_1
XFILLER_43_816 VPWR VGND sg13g2_decap_8
XFILLER_28_879 VPWR VGND sg13g2_decap_8
XFILLER_23_551 VPWR VGND sg13g2_decap_4
XFILLER_11_702 VPWR VGND sg13g2_fill_1
XFILLER_24_66 VPWR VGND sg13g2_decap_4
XFILLER_23_595 VPWR VGND sg13g2_fill_2
XFILLER_6_216 VPWR VGND sg13g2_fill_1
XFILLER_11_779 VPWR VGND sg13g2_fill_1
XFILLER_3_978 VPWR VGND sg13g2_decap_8
X_6136__312 VPWR VGND net312 sg13g2_tiehi
XFILLER_2_477 VPWR VGND sg13g2_fill_2
Xhold290 mydesign.accum\[78\] VPWR VGND net909 sg13g2_dlygate4sd3_1
XFILLER_19_824 VPWR VGND sg13g2_fill_1
XFILLER_37_109 VPWR VGND sg13g2_decap_8
XFILLER_46_621 VPWR VGND sg13g2_decap_8
XFILLER_18_323 VPWR VGND sg13g2_decap_4
XFILLER_45_142 VPWR VGND sg13g2_decap_8
XFILLER_46_698 VPWR VGND sg13g2_decap_8
XFILLER_45_164 VPWR VGND sg13g2_fill_2
X_3570_ VGND VPWR _0594_ _0595_ _0596_ net500 sg13g2_a21oi_1
XFILLER_6_783 VPWR VGND sg13g2_decap_4
X_5240_ VGND VPWR _2067_ _2068_ _2071_ _2052_ sg13g2_a21oi_1
X_5171_ VGND VPWR _2006_ _2007_ _2008_ _0397_ sg13g2_a21oi_1
X_4122_ VGND VPWR mydesign.pe_weights\[62\] _1046_ _1082_ mydesign.accum\[90\] sg13g2_a21oi_1
X_4053_ mydesign.pe_inputs\[55\] net428 mydesign.accum\[102\] _1025_ VPWR VGND sg13g2_nand3_1
XFILLER_49_492 VPWR VGND sg13g2_decap_8
XFILLER_49_470 VPWR VGND sg13g2_decap_4
XFILLER_37_643 VPWR VGND sg13g2_fill_2
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_2
XFILLER_37_676 VPWR VGND sg13g2_fill_1
XFILLER_40_819 VPWR VGND sg13g2_fill_2
X_4955_ net478 VPWR _1811_ VGND net589 net921 sg13g2_o21ai_1
X_3906_ mydesign.pe_inputs\[59\] _0804_ mydesign.accum\[110\] _0894_ VPWR VGND sg13g2_nand3_1
X_4886_ VGND VPWR net583 _1759_ _0243_ _1760_ sg13g2_a21oi_1
XFILLER_32_381 VPWR VGND sg13g2_fill_2
X_3837_ _0829_ _0812_ _0828_ VPWR VGND sg13g2_nand2_1
X_3768_ _0772_ VPWR _0113_ VGND net601 _0769_ sg13g2_o21ai_1
X_5507_ _2288_ VPWR _2309_ VGND _2277_ _2289_ sg13g2_o21ai_1
X_3699_ VGND VPWR net577 _0708_ _0107_ _0709_ sg13g2_a21oi_1
X_5438_ net635 VPWR _2246_ VGND mydesign.pe_inputs\[6\] net444 sg13g2_o21ai_1
XFILLER_0_915 VPWR VGND sg13g2_decap_8
X_5369_ _2184_ _2168_ _2182_ VPWR VGND sg13g2_xnor2_1
XFILLER_47_429 VPWR VGND sg13g2_fill_1
XFILLER_47_418 VPWR VGND sg13g2_decap_8
X_5890__373 VPWR VGND net373 sg13g2_tiehi
XFILLER_35_21 VPWR VGND sg13g2_decap_8
XFILLER_35_32 VPWR VGND sg13g2_fill_2
XFILLER_43_668 VPWR VGND sg13g2_fill_1
XFILLER_43_657 VPWR VGND sg13g2_fill_2
XFILLER_11_521 VPWR VGND sg13g2_fill_1
XFILLER_7_547 VPWR VGND sg13g2_decap_4
XFILLER_3_775 VPWR VGND sg13g2_fill_2
XFILLER_20_1003 VPWR VGND sg13g2_decap_8
XFILLER_47_985 VPWR VGND sg13g2_decap_8
XFILLER_46_451 VPWR VGND sg13g2_decap_4
XFILLER_15_882 VPWR VGND sg13g2_fill_1
X_4740_ net535 _1537_ mydesign.accum\[62\] _1632_ VPWR VGND sg13g2_nand3_1
X_4671_ _1567_ _1549_ _1565_ VPWR VGND sg13g2_xnor2_1
X_3622_ _0640_ mydesign.weights\[1\]\[16\] net495 VPWR VGND sg13g2_nand2_1
X_3553_ _0579_ _0512_ _0520_ VPWR VGND sg13g2_nand2_1
XFILLER_6_580 VPWR VGND sg13g2_fill_2
XFILLER_44_0 VPWR VGND sg13g2_decap_8
X_3484_ net621 VPWR _0518_ VGND net485 _0517_ sg13g2_o21ai_1
X_5223_ VPWR _2054_ _2053_ VGND sg13g2_inv_1
X_5154_ _1990_ VPWR _1993_ VGND _1973_ _1986_ sg13g2_o21ai_1
X_4105_ net808 _1046_ _1067_ VPWR VGND sg13g2_and2_1
XFILLER_38_930 VPWR VGND sg13g2_decap_8
X_5085_ _1928_ _1926_ _1927_ VPWR VGND sg13g2_nand2_1
X_4036_ _1009_ mydesign.pe_inputs\[55\] _0926_ VPWR VGND sg13g2_nand2_1
XFILLER_40_616 VPWR VGND sg13g2_fill_1
X_5987_ net182 VGND VPWR _0213_ mydesign.pe_inputs\[29\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_36_1021 VPWR VGND sg13g2_decap_8
X_4938_ _1793_ _1792_ _1795_ VPWR VGND sg13g2_xor2_1
X_4869_ _1745_ _1743_ _1744_ VPWR VGND sg13g2_nand2_1
XFILLER_21_874 VPWR VGND sg13g2_fill_2
XFILLER_21_885 VPWR VGND sg13g2_fill_2
XFILLER_0_756 VPWR VGND sg13g2_decap_4
XFILLER_48_727 VPWR VGND sg13g2_decap_8
XFILLER_0_767 VPWR VGND sg13g2_decap_4
XFILLER_0_789 VPWR VGND sg13g2_decap_8
XFILLER_47_237 VPWR VGND sg13g2_fill_1
XFILLER_29_930 VPWR VGND sg13g2_decap_8
XFILLER_44_911 VPWR VGND sg13g2_decap_8
XFILLER_16_602 VPWR VGND sg13g2_decap_8
XFILLER_44_988 VPWR VGND sg13g2_decap_8
XFILLER_15_145 VPWR VGND sg13g2_fill_1
XFILLER_31_616 VPWR VGND sg13g2_fill_1
XFILLER_43_498 VPWR VGND sg13g2_decap_4
XFILLER_30_137 VPWR VGND sg13g2_fill_2
XFILLER_8_801 VPWR VGND sg13g2_decap_4
XFILLER_39_738 VPWR VGND sg13g2_fill_1
XFILLER_47_782 VPWR VGND sg13g2_decap_8
X_5910_ net337 VGND VPWR _0136_ mydesign.pe_weights\[48\] clknet_leaf_44_clk sg13g2_dfrbpq_2
XFILLER_19_473 VPWR VGND sg13g2_decap_4
XFILLER_35_922 VPWR VGND sg13g2_decap_8
XFILLER_34_432 VPWR VGND sg13g2_fill_1
X_5841_ net87 VGND VPWR net408 mydesign.cp2\[2\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_22_605 VPWR VGND sg13g2_fill_1
XFILLER_35_999 VPWR VGND sg13g2_decap_8
XFILLER_22_627 VPWR VGND sg13g2_decap_8
X_5772_ _2515_ net674 _2511_ VPWR VGND sg13g2_nand2_1
X_4723_ _1614_ _1615_ _1616_ VPWR VGND sg13g2_and2_1
X_4654_ net815 _1521_ net686 _1551_ VPWR VGND sg13g2_nand3_1
X_3605_ _0627_ _0628_ _0094_ VPWR VGND sg13g2_nor2_1
X_4585_ VGND VPWR _1473_ _1476_ _1494_ _1492_ sg13g2_a21oi_1
X_3536_ _0562_ _0559_ _0563_ VPWR VGND sg13g2_xor2_1
X_5206_ VGND VPWR _2038_ _2037_ _2036_ sg13g2_or2_1
X_3467_ net554 mydesign.inputs\[0\]\[26\] _0503_ VPWR VGND sg13g2_nor2b_1
X_3398_ net517 mydesign.accum\[35\] _0445_ VPWR VGND sg13g2_nor2b_1
X_5137_ VGND VPWR _1976_ _1978_ _1960_ _1957_ sg13g2_a21oi_2
X_5068_ _1910_ _1907_ _1912_ VPWR VGND sg13g2_xor2_1
X_4019_ _0993_ _0991_ _0992_ VPWR VGND sg13g2_nand2_1
XFILLER_26_988 VPWR VGND sg13g2_decap_8
XFILLER_41_958 VPWR VGND sg13g2_decap_8
XFILLER_4_303 VPWR VGND sg13g2_fill_2
XFILLER_0_542 VPWR VGND sg13g2_fill_1
XFILLER_36_708 VPWR VGND sg13g2_fill_2
XFILLER_35_207 VPWR VGND sg13g2_decap_8
XFILLER_29_793 VPWR VGND sg13g2_decap_4
XFILLER_44_785 VPWR VGND sg13g2_decap_8
XFILLER_16_476 VPWR VGND sg13g2_fill_2
XFILLER_17_999 VPWR VGND sg13g2_decap_8
XFILLER_43_273 VPWR VGND sg13g2_fill_1
XFILLER_32_936 VPWR VGND sg13g2_decap_8
XFILLER_40_980 VPWR VGND sg13g2_decap_8
X_6105__236 VPWR VGND net236 sg13g2_tiehi
XFILLER_8_642 VPWR VGND sg13g2_decap_4
XFILLER_7_174 VPWR VGND sg13g2_fill_2
Xhold108 mydesign.weights\[0\]\[17\] VPWR VGND net727 sg13g2_dlygate4sd3_1
X_4370_ VGND VPWR mydesign.pe_weights\[53\] net534 _1299_ mydesign.accum\[73\] sg13g2_a21oi_1
X_5940__277 VPWR VGND net277 sg13g2_tiehi
Xhold119 mydesign.inputs\[0\]\[27\] VPWR VGND net738 sg13g2_dlygate4sd3_1
X_3321_ _0376_ VPWR _0380_ VGND _2599_ _2656_ sg13g2_o21ai_1
X_3252_ net791 _2669_ _2659_ _0023_ VPWR VGND sg13g2_mux2_1
XFILLER_3_391 VPWR VGND sg13g2_decap_8
X_6040_ net298 VGND VPWR _0266_ mydesign.accum\[46\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_3183_ net1044 net842 _2619_ VPWR VGND sg13g2_nor2_2
XFILLER_27_708 VPWR VGND sg13g2_fill_1
XFILLER_35_774 VPWR VGND sg13g2_decap_8
X_5824_ net118 VGND VPWR _0050_ mydesign.inputs\[0\]\[17\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5755_ VGND VPWR _1771_ _2505_ _0365_ net824 sg13g2_a21oi_1
X_5686_ _2468_ net623 net430 VPWR VGND sg13g2_nand2_1
XFILLER_30_490 VPWR VGND sg13g2_fill_1
X_4706_ _1600_ _1598_ _1599_ VPWR VGND sg13g2_nand2_1
X_4637_ net623 VPWR _1539_ VGND net891 net439 sg13g2_o21ai_1
X_6119__84 VPWR VGND net84 sg13g2_tiehi
X_5802__148 VPWR VGND net148 sg13g2_tiehi
X_4568_ net473 VPWR _1478_ VGND net574 net841 sg13g2_o21ai_1
X_4499_ VGND VPWR net690 _1411_ _0204_ _1412_ sg13g2_a21oi_1
X_3519_ _0547_ _0546_ _0530_ VPWR VGND sg13g2_nand2b_1
XFILLER_17_218 VPWR VGND sg13g2_fill_2
XFILLER_14_914 VPWR VGND sg13g2_fill_1
XFILLER_43_65 VPWR VGND sg13g2_fill_1
XFILLER_9_417 VPWR VGND sg13g2_fill_2
XFILLER_40_265 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_20_clk clknet_3_3__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_5_612 VPWR VGND sg13g2_decap_4
XFILLER_4_133 VPWR VGND sg13g2_fill_1
X_6125__32 VPWR VGND net32 sg13g2_tiehi
XFILLER_1_840 VPWR VGND sg13g2_fill_1
XFILLER_1_851 VPWR VGND sg13g2_fill_1
XFILLER_49_811 VPWR VGND sg13g2_decap_8
XFILLER_0_361 VPWR VGND sg13g2_decap_8
XFILLER_0_383 VPWR VGND sg13g2_fill_2
XFILLER_49_888 VPWR VGND sg13g2_decap_8
XFILLER_16_240 VPWR VGND sg13g2_fill_2
XFILLER_17_752 VPWR VGND sg13g2_fill_2
XFILLER_32_722 VPWR VGND sg13g2_fill_1
XFILLER_16_295 VPWR VGND sg13g2_fill_2
X_3870_ mydesign.pe_inputs\[57\] _0804_ mydesign.accum\[108\] _0860_ VPWR VGND sg13g2_nand3_1
XFILLER_13_980 VPWR VGND sg13g2_decap_8
X_5540_ _2322_ _2321_ _2338_ _2340_ VPWR VGND sg13g2_a21o_1
Xclkbuf_leaf_11_clk clknet_3_2__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
XFILLER_9_984 VPWR VGND sg13g2_decap_8
X_5471_ VGND VPWR net588 _2273_ _0314_ _2274_ sg13g2_a21oi_1
X_4422_ mydesign.pe_inputs\[41\] net538 mydesign.accum\[76\] _1348_ VPWR VGND sg13g2_a21o_1
X_4353_ VGND VPWR _2562_ net433 _0181_ _1289_ sg13g2_a21oi_1
X_4284_ _1226_ _1209_ _1227_ VPWR VGND sg13g2_nor2b_1
Xfanout429 _2692_ net429 VPWR VGND sg13g2_buf_8
X_3304_ net605 _2656_ net1064 _2692_ VPWR VGND sg13g2_nand3_1
X_6023_ net370 VGND VPWR net860 mydesign.weights\[3\]\[9\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3235_ _2655_ net614 _2618_ VPWR VGND sg13g2_nand2_2
XFILLER_39_376 VPWR VGND sg13g2_fill_1
X_3166_ _2606_ net1106 VPWR VGND mydesign.load_counter\[0\] sg13g2_nand2b_2
X_3097_ VPWR _2538_ net1031 VGND sg13g2_inv_1
X_3999_ VGND VPWR _0971_ _0972_ _0974_ _0951_ sg13g2_a21oi_1
X_5807_ net139 VGND VPWR _0033_ mydesign.inputs\[2\]\[16\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_13_46 VPWR VGND sg13g2_decap_8
X_5738_ _2498_ net694 _2495_ VPWR VGND sg13g2_nand2_1
X_5669_ VGND VPWR mydesign.accum\[6\] _2445_ _2456_ _2447_ sg13g2_a21oi_1
Xhold472 mydesign.pe_weights\[48\] VPWR VGND net1091 sg13g2_dlygate4sd3_1
Xhold450 net9 VPWR VGND net1069 sg13g2_dlygate4sd3_1
Xhold461 net13 VPWR VGND net1080 sg13g2_dlygate4sd3_1
X_5919__319 VPWR VGND net319 sg13g2_tiehi
Xhold483 mydesign.pe_inputs\[60\] VPWR VGND net1102 sg13g2_dlygate4sd3_1
XFILLER_46_803 VPWR VGND sg13g2_decap_8
XFILLER_18_516 VPWR VGND sg13g2_fill_1
XFILLER_14_755 VPWR VGND sg13g2_fill_2
XFILLER_26_593 VPWR VGND sg13g2_decap_4
Xclkload17 clknet_leaf_27_clk clkload17/X VPWR VGND sg13g2_buf_8
XFILLER_6_965 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_23_1001 VPWR VGND sg13g2_decap_8
XFILLER_49_685 VPWR VGND sg13g2_decap_8
XFILLER_37_825 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_24_519 VPWR VGND sg13g2_decap_4
XFILLER_45_891 VPWR VGND sg13g2_decap_8
X_4971_ _1826_ _1802_ _1824_ VPWR VGND sg13g2_xnor2_1
X_3922_ net472 VPWR _0909_ VGND net578 net835 sg13g2_o21ai_1
X_3853_ _0844_ _0820_ _0842_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_574 VPWR VGND sg13g2_fill_2
XFILLER_20_736 VPWR VGND sg13g2_fill_1
XFILLER_9_770 VPWR VGND sg13g2_fill_1
X_3784_ net459 VPWR _0782_ VGND net552 mydesign.weights\[2\]\[8\] sg13g2_o21ai_1
XFILLER_20_769 VPWR VGND sg13g2_fill_2
X_5523_ _2303_ VPWR _2324_ VGND _2296_ _2304_ sg13g2_o21ai_1
X_5454_ net477 VPWR _2259_ VGND net588 net928 sg13g2_o21ai_1
X_5385_ _2176_ _2178_ _2197_ _2199_ VPWR VGND sg13g2_or3_1
X_4405_ _1310_ _1331_ _1332_ VPWR VGND sg13g2_nor2b_1
X_4336_ _1258_ _1275_ _1257_ _1276_ VPWR VGND sg13g2_nand3_1
X_4267_ _1201_ VPWR _1210_ VGND _1194_ _1202_ sg13g2_o21ai_1
X_4198_ VGND VPWR _1139_ _1153_ _1155_ net500 sg13g2_a21oi_1
X_3218_ _2644_ VPWR _0014_ VGND net602 _2641_ sg13g2_o21ai_1
X_6006_ net70 VGND VPWR net1014 mydesign.pe_weights\[24\] clknet_leaf_29_clk sg13g2_dfrbpq_2
XFILLER_39_184 VPWR VGND sg13g2_fill_2
XFILLER_39_162 VPWR VGND sg13g2_decap_4
X_3149_ VPWR _2590_ net623 VGND sg13g2_inv_1
XFILLER_27_357 VPWR VGND sg13g2_decap_8
XFILLER_24_12 VPWR VGND sg13g2_fill_1
X_6025__362 VPWR VGND net362 sg13g2_tiehi
XFILLER_10_257 VPWR VGND sg13g2_fill_2
XFILLER_10_268 VPWR VGND sg13g2_fill_2
X_6095__316 VPWR VGND net316 sg13g2_tiehi
XFILLER_2_401 VPWR VGND sg13g2_fill_2
XFILLER_3_957 VPWR VGND sg13g2_decap_8
Xhold280 mydesign.pe_inputs\[41\] VPWR VGND net899 sg13g2_dlygate4sd3_1
XFILLER_49_64 VPWR VGND sg13g2_fill_1
Xhold291 mydesign.pe_weights\[52\] VPWR VGND net910 sg13g2_dlygate4sd3_1
XFILLER_46_600 VPWR VGND sg13g2_decap_8
XFILLER_1_38 VPWR VGND sg13g2_fill_2
XFILLER_46_677 VPWR VGND sg13g2_decap_8
XFILLER_5_261 VPWR VGND sg13g2_decap_8
X_5170_ _2007_ net549 mydesign.inputs\[3\]\[5\] VPWR VGND sg13g2_nand2_1
X_4121_ _1081_ mydesign.accum\[90\] mydesign.pe_weights\[62\] _1046_ VPWR VGND sg13g2_and3_2
X_6072__168 VPWR VGND net168 sg13g2_tiehi
X_4052_ VGND VPWR mydesign.pe_inputs\[55\] net428 _1024_ mydesign.accum\[102\] sg13g2_a21oi_1
X_6113__176 VPWR VGND net176 sg13g2_tiehi
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_2
XFILLER_37_666 VPWR VGND sg13g2_fill_2
XFILLER_25_817 VPWR VGND sg13g2_fill_2
XFILLER_40_809 VPWR VGND sg13g2_fill_2
X_4954_ _1810_ _1794_ _1809_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_338 VPWR VGND sg13g2_decap_4
X_3905_ VGND VPWR mydesign.pe_inputs\[59\] _0804_ _0893_ mydesign.accum\[110\] sg13g2_a21oi_1
X_4885_ net479 VPWR _1760_ VGND net590 net912 sg13g2_o21ai_1
X_3836_ _0828_ _0818_ _0826_ VPWR VGND sg13g2_xnor2_1
X_3767_ _0772_ net672 _0770_ VPWR VGND sg13g2_nand2_1
XFILLER_20_588 VPWR VGND sg13g2_fill_1
X_5506_ _2306_ _2307_ _2308_ VPWR VGND sg13g2_and2_1
X_3698_ net470 VPWR _0709_ VGND net577 net936 sg13g2_o21ai_1
X_5437_ VGND VPWR _2523_ net444 _0309_ _2245_ sg13g2_a21oi_1
X_5368_ _2168_ _2182_ _2183_ VPWR VGND sg13g2_and2_1
XFILLER_48_909 VPWR VGND sg13g2_decap_8
X_4319_ _1258_ _1257_ _1260_ VPWR VGND sg13g2_xor2_1
X_5299_ _2125_ net837 _2126_ VPWR VGND sg13g2_xor2_1
XFILLER_19_56 VPWR VGND sg13g2_decap_4
XFILLER_16_806 VPWR VGND sg13g2_fill_2
XFILLER_27_143 VPWR VGND sg13g2_decap_4
XFILLER_42_102 VPWR VGND sg13g2_fill_1
XFILLER_42_124 VPWR VGND sg13g2_decap_8
XFILLER_42_113 VPWR VGND sg13g2_fill_1
XFILLER_42_157 VPWR VGND sg13g2_decap_8
XFILLER_24_883 VPWR VGND sg13g2_decap_8
XFILLER_11_533 VPWR VGND sg13g2_decap_8
XFILLER_13_1022 VPWR VGND sg13g2_decap_8
XFILLER_3_721 VPWR VGND sg13g2_decap_4
XFILLER_4_0 VPWR VGND sg13g2_fill_2
Xfanout590 net591 net590 VPWR VGND sg13g2_buf_8
XFILLER_47_964 VPWR VGND sg13g2_decap_8
XFILLER_18_121 VPWR VGND sg13g2_fill_2
XFILLER_33_135 VPWR VGND sg13g2_decap_4
XFILLER_33_168 VPWR VGND sg13g2_fill_2
XFILLER_41_190 VPWR VGND sg13g2_decap_8
XFILLER_14_393 VPWR VGND sg13g2_fill_2
X_6004__78 VPWR VGND net78 sg13g2_tiehi
XFILLER_30_842 VPWR VGND sg13g2_fill_1
X_4670_ _1566_ _1549_ _1565_ VPWR VGND sg13g2_nand2_1
X_3621_ net556 _0397_ _0639_ VPWR VGND sg13g2_nor2_2
X_3552_ _0578_ _0564_ _0566_ VPWR VGND sg13g2_nand2_1
X_3483_ VGND VPWR net543 _0517_ _0516_ _0515_ sg13g2_a21oi_2
X_5222_ _2053_ mydesign.pe_weights\[28\] _2020_ VPWR VGND sg13g2_nand2_1
X_5153_ VGND VPWR net575 _1991_ _0278_ _1992_ sg13g2_a21oi_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
X_4104_ VGND VPWR _2575_ net437 _0155_ _1066_ sg13g2_a21oi_1
X_5084_ mydesign.pe_inputs\[21\] mydesign.pe_weights\[34\] mydesign.accum\[35\] _1927_
+ VPWR VGND sg13g2_a21o_1
X_5950__257 VPWR VGND net257 sg13g2_tiehi
X_4035_ _0995_ VPWR _1008_ VGND _0988_ _0996_ sg13g2_o21ai_1
XFILLER_38_986 VPWR VGND sg13g2_decap_8
XFILLER_25_669 VPWR VGND sg13g2_decap_8
X_5986_ net185 VGND VPWR _0212_ mydesign.pe_inputs\[28\] clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_36_1000 VPWR VGND sg13g2_decap_8
X_4937_ mydesign.pe_weights\[36\] net528 net664 _1794_ VPWR VGND _1792_ sg13g2_nand4_1
X_4868_ mydesign.pe_inputs\[31\] mydesign.pe_weights\[43\] mydesign.accum\[54\] _1744_
+ VPWR VGND sg13g2_a21o_1
XFILLER_32_190 VPWR VGND sg13g2_fill_1
X_3819_ _0810_ _0811_ _0812_ VPWR VGND sg13g2_nor2_1
XFILLER_21_13 VPWR VGND sg13g2_decap_8
X_4799_ _1679_ _1661_ _1678_ VPWR VGND sg13g2_nand2_1
XFILLER_48_706 VPWR VGND sg13g2_decap_8
XFILLER_43_1026 VPWR VGND sg13g2_fill_2
XFILLER_29_986 VPWR VGND sg13g2_decap_8
XFILLER_46_87 VPWR VGND sg13g2_fill_2
XFILLER_44_967 VPWR VGND sg13g2_decap_8
XFILLER_28_496 VPWR VGND sg13g2_decap_4
XFILLER_43_455 VPWR VGND sg13g2_fill_1
XFILLER_24_680 VPWR VGND sg13g2_fill_1
XFILLER_12_842 VPWR VGND sg13g2_fill_2
XFILLER_7_334 VPWR VGND sg13g2_fill_1
XFILLER_30_7 VPWR VGND sg13g2_fill_1
XFILLER_47_761 VPWR VGND sg13g2_decap_8
XFILLER_19_463 VPWR VGND sg13g2_fill_2
XFILLER_35_901 VPWR VGND sg13g2_decap_8
XFILLER_34_422 VPWR VGND sg13g2_decap_4
X_5840_ net89 VGND VPWR _0066_ mydesign.cp2\[1\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_35_978 VPWR VGND sg13g2_decap_8
X_5771_ _2514_ VPWR _0374_ VGND net600 _2511_ sg13g2_o21ai_1
X_5828__113 VPWR VGND net113 sg13g2_tiehi
XFILLER_30_650 VPWR VGND sg13g2_fill_1
X_4722_ _2548_ VPWR _1615_ VGND _2549_ _1531_ sg13g2_o21ai_1
X_4653_ _1548_ _1547_ _1550_ VPWR VGND sg13g2_xor2_1
X_3604_ net468 VPWR _0628_ VGND net558 net1062 sg13g2_o21ai_1
X_4584_ _1493_ _1473_ _1476_ _1492_ VPWR VGND sg13g2_and3_1
X_3535_ _0560_ mydesign.accum\[123\] _0562_ VPWR VGND sg13g2_xor2_1
X_3466_ net609 _0502_ _0081_ VPWR VGND sg13g2_nor2_1
X_5205_ VGND VPWR mydesign.pe_weights\[30\] _2004_ _2037_ mydesign.accum\[26\] sg13g2_a21oi_1
X_3397_ mydesign.accum\[99\] mydesign.accum\[67\] net512 _0444_ VPWR VGND sg13g2_mux2_1
X_6091__352 VPWR VGND net352 sg13g2_tiehi
X_5136_ _1977_ _1957_ _1960_ _1976_ VPWR VGND sg13g2_and3_1
XFILLER_45_709 VPWR VGND sg13g2_decap_8
XFILLER_38_750 VPWR VGND sg13g2_fill_2
X_5067_ _1907_ _1910_ _1911_ VPWR VGND sg13g2_nor2_1
XFILLER_38_783 VPWR VGND sg13g2_fill_1
XFILLER_38_772 VPWR VGND sg13g2_fill_2
X_4018_ _0933_ mydesign.pe_inputs\[53\] mydesign.accum\[100\] _0992_ VPWR VGND sg13g2_a21o_1
XFILLER_37_260 VPWR VGND sg13g2_fill_2
XFILLER_25_411 VPWR VGND sg13g2_decap_4
XFILLER_26_967 VPWR VGND sg13g2_decap_8
XFILLER_16_68 VPWR VGND sg13g2_fill_1
XFILLER_25_444 VPWR VGND sg13g2_fill_2
XFILLER_41_937 VPWR VGND sg13g2_decap_8
X_5969_ net219 VGND VPWR _0195_ mydesign.accum\[79\] clknet_leaf_31_clk sg13g2_dfrbpq_1
XFILLER_0_521 VPWR VGND sg13g2_decap_8
XFILLER_48_547 VPWR VGND sg13g2_decap_4
XFILLER_44_764 VPWR VGND sg13g2_decap_8
XFILLER_43_252 VPWR VGND sg13g2_fill_2
XFILLER_16_455 VPWR VGND sg13g2_fill_1
XFILLER_17_978 VPWR VGND sg13g2_decap_8
XFILLER_32_915 VPWR VGND sg13g2_decap_8
XFILLER_31_458 VPWR VGND sg13g2_fill_1
XFILLER_12_661 VPWR VGND sg13g2_fill_1
XFILLER_11_182 VPWR VGND sg13g2_fill_1
XFILLER_8_687 VPWR VGND sg13g2_fill_1
X_5905__343 VPWR VGND net343 sg13g2_tiehi
Xhold109 mydesign.inputs\[0\]\[26\] VPWR VGND net728 sg13g2_dlygate4sd3_1
X_3320_ VGND VPWR _0378_ _0379_ _0058_ net607 sg13g2_a21oi_1
X_3251_ net3 _2666_ _2669_ VPWR VGND sg13g2_and2_1
X_3182_ _2618_ _2591_ net5 VPWR VGND sg13g2_nand2_2
XFILLER_39_558 VPWR VGND sg13g2_fill_2
XFILLER_14_2 VPWR VGND sg13g2_fill_1
XFILLER_34_230 VPWR VGND sg13g2_fill_2
X_5823_ net119 VGND VPWR _0049_ mydesign.inputs\[0\]\[16\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_23_959 VPWR VGND sg13g2_decap_8
X_5754_ net612 VPWR _2507_ VGND net823 _2505_ sg13g2_o21ai_1
X_5685_ net608 _2698_ _2467_ VPWR VGND sg13g2_nor2_1
XFILLER_31_992 VPWR VGND sg13g2_decap_8
X_4705_ _1527_ net535 mydesign.accum\[60\] _1599_ VPWR VGND sg13g2_a21o_1
XFILLER_8_80 VPWR VGND sg13g2_fill_1
X_4636_ VGND VPWR _2545_ net493 _0215_ _1538_ sg13g2_a21oi_1
X_4567_ VGND VPWR _1475_ _1476_ _1477_ net501 sg13g2_a21oi_1
X_4498_ net473 VPWR _1412_ VGND net690 _1411_ sg13g2_o21ai_1
X_3518_ _0544_ _0543_ _0546_ VPWR VGND sg13g2_xor2_1
X_3449_ _2639_ _2683_ _0491_ VPWR VGND sg13g2_nor2_1
X_5119_ VGND VPWR _1959_ _1960_ _1961_ net503 sg13g2_a21oi_1
XFILLER_45_528 VPWR VGND sg13g2_fill_1
XFILLER_45_517 VPWR VGND sg13g2_fill_1
XFILLER_45_506 VPWR VGND sg13g2_fill_2
X_6099_ net284 VGND VPWR net1058 mydesign.accum\[1\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_26_731 VPWR VGND sg13g2_fill_1
XFILLER_25_241 VPWR VGND sg13g2_decap_8
XFILLER_40_244 VPWR VGND sg13g2_fill_2
XFILLER_13_447 VPWR VGND sg13g2_fill_1
XFILLER_49_1021 VPWR VGND sg13g2_decap_8
XFILLER_48_300 VPWR VGND sg13g2_decap_4
XFILLER_1_874 VPWR VGND sg13g2_fill_1
XFILLER_49_867 VPWR VGND sg13g2_decap_8
XFILLER_48_355 VPWR VGND sg13g2_fill_1
XFILLER_16_230 VPWR VGND sg13g2_fill_1
XFILLER_31_255 VPWR VGND sg13g2_fill_2
XFILLER_31_266 VPWR VGND sg13g2_fill_1
XFILLER_9_963 VPWR VGND sg13g2_decap_8
X_5470_ net477 VPWR _2274_ VGND net588 net1038 sg13g2_o21ai_1
X_4421_ net538 mydesign.pe_inputs\[41\] mydesign.accum\[76\] _1347_ VPWR VGND sg13g2_nand3_1
X_4352_ net628 VPWR _1289_ VGND net966 net434 sg13g2_o21ai_1
X_4283_ _1226_ _1210_ _1224_ VPWR VGND sg13g2_xnor2_1
X_3303_ net801 _2670_ _2691_ _0052_ VPWR VGND sg13g2_mux2_1
X_6022_ net378 VGND VPWR net846 mydesign.weights\[3\]\[8\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3234_ _2654_ VPWR _0020_ VGND net598 _2649_ sg13g2_o21ai_1
X_3165_ _2605_ net614 net610 VPWR VGND sg13g2_nand2_2
X_3096_ VPWR _2537_ net974 VGND sg13g2_inv_1
XFILLER_35_561 VPWR VGND sg13g2_fill_2
X_3998_ _0973_ _0951_ _0971_ _0972_ VPWR VGND sg13g2_and3_1
X_5806_ net141 VGND VPWR _0032_ mydesign.weights\[2\]\[15\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_22_244 VPWR VGND sg13g2_decap_8
XFILLER_22_266 VPWR VGND sg13g2_decap_8
X_5737_ _2497_ VPWR _0357_ VGND net602 _2495_ sg13g2_o21ai_1
X_5668_ VGND VPWR net587 _2454_ _0330_ _2455_ sg13g2_a21oi_1
X_5599_ _2377_ VPWR _2390_ VGND _2375_ _2378_ sg13g2_o21ai_1
XFILLER_2_605 VPWR VGND sg13g2_fill_2
X_4619_ _1524_ _0392_ _1523_ VPWR VGND sg13g2_nand2_1
Xhold451 _0069_ VPWR VGND net1070 sg13g2_dlygate4sd3_1
Xhold462 net8 VPWR VGND net1081 sg13g2_dlygate4sd3_1
Xhold440 mydesign.pe_inputs\[63\] VPWR VGND net1059 sg13g2_dlygate4sd3_1
Xhold484 mydesign.out\[3\] VPWR VGND net1103 sg13g2_dlygate4sd3_1
Xhold473 mydesign.pe_weights\[55\] VPWR VGND net1092 sg13g2_dlygate4sd3_1
X_5776__181 VPWR VGND net181 sg13g2_tiehi
XFILLER_46_859 VPWR VGND sg13g2_decap_8
XFILLER_14_745 VPWR VGND sg13g2_decap_4
XFILLER_13_266 VPWR VGND sg13g2_fill_1
XFILLER_13_299 VPWR VGND sg13g2_fill_1
XFILLER_10_984 VPWR VGND sg13g2_decap_8
Xclkload18 VPWR clkload18/Y clknet_leaf_33_clk VGND sg13g2_inv_1
XFILLER_0_181 VPWR VGND sg13g2_fill_2
XFILLER_49_664 VPWR VGND sg13g2_decap_8
XFILLER_45_870 VPWR VGND sg13g2_decap_8
X_4970_ _1825_ _1802_ _1824_ VPWR VGND sg13g2_nand2_1
XFILLER_44_380 VPWR VGND sg13g2_fill_1
X_3921_ _0908_ _0904_ _0907_ VPWR VGND sg13g2_xnor2_1
X_3852_ VPWR _0843_ _0842_ VGND sg13g2_inv_1
X_3783_ net497 mydesign.weights\[2\]\[4\] _0781_ VPWR VGND sg13g2_nor2_1
X_5522_ _2322_ _2321_ _2323_ VPWR VGND sg13g2_xor2_1
X_5453_ _2256_ _2255_ _2258_ VPWR VGND sg13g2_xor2_1
X_5384_ _2197_ VPWR _2198_ VGND _2176_ _2178_ sg13g2_o21ai_1
X_4404_ _1330_ _1327_ _1331_ VPWR VGND sg13g2_xor2_1
X_4335_ _1273_ _1274_ _1275_ VPWR VGND sg13g2_and2_1
X_4266_ _1205_ VPWR _1209_ VGND _1191_ _1206_ sg13g2_o21ai_1
X_4197_ VGND VPWR _1154_ _1153_ _1139_ sg13g2_or2_1
X_3217_ _2644_ net420 _2642_ VPWR VGND sg13g2_nand2_1
X_6005_ net74 VGND VPWR net888 mydesign.pe_inputs\[27\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_3148_ VPWR _2589_ mydesign.weights\[2\]\[16\] VGND sg13g2_inv_1
X_3079_ _2520_ net1 VPWR VGND sg13g2_inv_2
XFILLER_11_726 VPWR VGND sg13g2_fill_2
XFILLER_23_586 VPWR VGND sg13g2_fill_1
X_5960__237 VPWR VGND net237 sg13g2_tiehi
XFILLER_3_903 VPWR VGND sg13g2_decap_4
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_46_1013 VPWR VGND sg13g2_decap_8
Xhold270 mydesign.accum\[39\] VPWR VGND net889 sg13g2_dlygate4sd3_1
XFILLER_49_54 VPWR VGND sg13g2_fill_1
XFILLER_49_43 VPWR VGND sg13g2_decap_8
Xhold292 mydesign.accum\[83\] VPWR VGND net911 sg13g2_dlygate4sd3_1
Xhold281 mydesign.accum\[50\] VPWR VGND net900 sg13g2_dlygate4sd3_1
XFILLER_46_656 VPWR VGND sg13g2_decap_8
XFILLER_45_166 VPWR VGND sg13g2_fill_1
XFILLER_27_881 VPWR VGND sg13g2_fill_1
XFILLER_45_199 VPWR VGND sg13g2_fill_1
XFILLER_42_884 VPWR VGND sg13g2_decap_8
X_6065__198 VPWR VGND net198 sg13g2_tiehi
X_4120_ _1080_ mydesign.pe_weights\[60\] _1056_ VPWR VGND sg13g2_nand2_1
X_4051_ _1022_ VPWR _1023_ VGND _1004_ _1019_ sg13g2_o21ai_1
XFILLER_49_461 VPWR VGND sg13g2_decap_4
X_5845__79 VPWR VGND net79 sg13g2_tiehi
Xinput5 ui_in[5] net5 VPWR VGND sg13g2_buf_2
XFILLER_37_645 VPWR VGND sg13g2_fill_1
X_4953_ _1809_ _1790_ _1807_ VPWR VGND sg13g2_xnor2_1
X_3904_ _0888_ VPWR _0892_ VGND _0876_ _0889_ sg13g2_o21ai_1
XFILLER_32_350 VPWR VGND sg13g2_decap_4
X_4884_ _1759_ _1755_ _1758_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_383 VPWR VGND sg13g2_fill_1
X_3835_ _0827_ _0826_ _0818_ VPWR VGND sg13g2_nand2b_1
X_3766_ _0771_ VPWR _0112_ VGND net603 _0769_ sg13g2_o21ai_1
X_5505_ _2284_ _2286_ _2305_ _2307_ VPWR VGND sg13g2_or3_1
X_5436_ net635 VPWR _2245_ VGND mydesign.pe_inputs\[5\] net444 sg13g2_o21ai_1
X_3697_ _0708_ _0687_ _0707_ VPWR VGND sg13g2_xnor2_1
X_5367_ _2181_ _2169_ _2182_ VPWR VGND sg13g2_xor2_1
X_4318_ _1259_ _1257_ _1258_ VPWR VGND sg13g2_nand2_1
X_5298_ _2112_ VPWR _2125_ VGND _2111_ _2115_ sg13g2_o21ai_1
X_4249_ VGND VPWR net570 _1192_ _0173_ _1193_ sg13g2_a21oi_1
XFILLER_27_100 VPWR VGND sg13g2_fill_2
XFILLER_28_623 VPWR VGND sg13g2_decap_4
XFILLER_27_122 VPWR VGND sg13g2_decap_8
XFILLER_13_1001 VPWR VGND sg13g2_decap_8
XFILLER_7_516 VPWR VGND sg13g2_decap_4
XFILLER_3_744 VPWR VGND sg13g2_fill_1
X_6071__180 VPWR VGND net180 sg13g2_tiehi
Xfanout580 net581 net580 VPWR VGND sg13g2_buf_2
Xfanout591 net593 net591 VPWR VGND sg13g2_buf_8
XFILLER_47_943 VPWR VGND sg13g2_decap_8
XFILLER_46_420 VPWR VGND sg13g2_decap_8
XFILLER_34_604 VPWR VGND sg13g2_decap_8
XFILLER_21_309 VPWR VGND sg13g2_decap_4
X_3620_ VGND VPWR _2580_ net490 _0099_ _0638_ sg13g2_a21oi_1
X_3551_ _0576_ _0577_ _0091_ VPWR VGND sg13g2_nor2_1
X_3482_ _0516_ _0394_ mydesign.weights\[0\]\[12\] net496 mydesign.weights\[0\]\[16\]
+ VPWR VGND sg13g2_a22oi_1
X_5221_ _2052_ _2042_ _2044_ VPWR VGND sg13g2_nand2_1
X_5152_ net474 VPWR _1992_ VGND net575 net826 sg13g2_o21ai_1
X_4103_ net624 VPWR _1066_ VGND net927 net436 sg13g2_o21ai_1
X_5083_ mydesign.pe_weights\[34\] mydesign.pe_inputs\[21\] mydesign.accum\[35\] _1926_
+ VPWR VGND sg13g2_nand3_1
XFILLER_38_965 VPWR VGND sg13g2_decap_8
X_4034_ _1007_ _1001_ _1004_ VPWR VGND sg13g2_nand2_1
XFILLER_40_607 VPWR VGND sg13g2_decap_8
X_5985_ net187 VGND VPWR _0211_ mydesign.accum\[71\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_4936_ net943 net528 net664 _1793_ VPWR VGND sg13g2_nand3_1
X_4867_ net533 mydesign.pe_inputs\[31\] mydesign.accum\[54\] _1743_ VPWR VGND sg13g2_nand3_1
XFILLER_20_331 VPWR VGND sg13g2_decap_8
XFILLER_21_865 VPWR VGND sg13g2_fill_1
X_3818_ _0811_ mydesign.pe_inputs\[57\] _0783_ VPWR VGND sg13g2_nand2_1
XFILLER_20_353 VPWR VGND sg13g2_decap_8
XFILLER_21_876 VPWR VGND sg13g2_fill_1
XFILLER_21_887 VPWR VGND sg13g2_fill_1
X_4798_ _1678_ _1668_ _1677_ VPWR VGND sg13g2_xnor2_1
X_3749_ _0723_ _0743_ _0757_ VPWR VGND sg13g2_nor2_1
X_5419_ _2231_ _2230_ _2229_ VPWR VGND sg13g2_nand2b_1
XFILLER_43_1005 VPWR VGND sg13g2_decap_8
XFILLER_0_725 VPWR VGND sg13g2_decap_8
XFILLER_28_431 VPWR VGND sg13g2_fill_1
XFILLER_29_965 VPWR VGND sg13g2_decap_8
XFILLER_44_946 VPWR VGND sg13g2_decap_8
XFILLER_16_648 VPWR VGND sg13g2_fill_2
XFILLER_8_825 VPWR VGND sg13g2_fill_2
XFILLER_11_375 VPWR VGND sg13g2_fill_1
XFILLER_8_869 VPWR VGND sg13g2_fill_1
XFILLER_7_379 VPWR VGND sg13g2_fill_2
XFILLER_7_368 VPWR VGND sg13g2_decap_8
X_5897__359 VPWR VGND net359 sg13g2_tiehi
XFILLER_47_740 VPWR VGND sg13g2_decap_8
XFILLER_35_957 VPWR VGND sg13g2_decap_8
X_5770_ _2514_ net737 _2511_ VPWR VGND sg13g2_nand2_1
XFILLER_30_640 VPWR VGND sg13g2_fill_2
X_4721_ net535 mydesign.accum\[61\] _1614_ VPWR VGND _1531_ sg13g2_nand3b_1
X_4652_ _1547_ _1548_ _1549_ VPWR VGND sg13g2_nor2_1
X_3603_ VGND VPWR _0625_ _0626_ _0627_ net500 sg13g2_a21oi_1
X_4583_ _1490_ _1469_ _1492_ VPWR VGND sg13g2_xor2_1
X_3534_ _0498_ _0526_ mydesign.accum\[123\] _0561_ VPWR VGND sg13g2_nand3_1
X_3465_ _0502_ _0499_ _0501_ net484 net1071 VPWR VGND sg13g2_a22oi_1
X_5204_ _2036_ mydesign.accum\[26\] mydesign.pe_weights\[30\] _2004_ VPWR VGND sg13g2_and3_1
X_3396_ net513 mydesign.accum\[107\] mydesign.accum\[75\] mydesign.accum\[43\] mydesign.accum\[11\]
+ net506 _0443_ VPWR VGND sg13g2_mux4_1
X_5135_ _1976_ _1953_ _1974_ VPWR VGND sg13g2_xnor2_1
X_5066_ _1910_ _1908_ _1909_ VPWR VGND sg13g2_nand2_1
X_4017_ mydesign.pe_inputs\[53\] net428 mydesign.accum\[100\] _0991_ VPWR VGND sg13g2_nand3_1
X_6082__52 VPWR VGND net52 sg13g2_tiehi
XFILLER_26_946 VPWR VGND sg13g2_decap_8
XFILLER_37_272 VPWR VGND sg13g2_fill_2
XFILLER_37_294 VPWR VGND sg13g2_decap_8
XFILLER_41_916 VPWR VGND sg13g2_decap_8
X_5968_ net221 VGND VPWR _0194_ mydesign.accum\[78\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_4919_ net635 VPWR _1781_ VGND net1043 net444 sg13g2_o21ai_1
X_5899_ net355 VGND VPWR net917 mydesign.accum\[105\] clknet_leaf_41_clk sg13g2_dfrbpq_2
XFILLER_21_673 VPWR VGND sg13g2_decap_8
XFILLER_10_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_588 VPWR VGND sg13g2_decap_4
XFILLER_17_902 VPWR VGND sg13g2_fill_2
XFILLER_17_957 VPWR VGND sg13g2_decap_8
XFILLER_44_743 VPWR VGND sg13g2_decap_8
XFILLER_43_264 VPWR VGND sg13g2_decap_8
XFILLER_7_121 VPWR VGND sg13g2_fill_1
XFILLER_4_861 VPWR VGND sg13g2_fill_1
X_3250_ net799 _2668_ _2659_ _0022_ VPWR VGND sg13g2_mux2_1
X_3181_ net610 net5 _2617_ VPWR VGND sg13g2_nor2b_2
XFILLER_21_4 VPWR VGND sg13g2_decap_4
XFILLER_34_242 VPWR VGND sg13g2_decap_8
X_5822_ net120 VGND VPWR _0048_ mydesign.inputs\[0\]\[15\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_22_415 VPWR VGND sg13g2_fill_1
XFILLER_34_253 VPWR VGND sg13g2_fill_1
X_5753_ VGND VPWR _1769_ _2505_ _0364_ net986 sg13g2_a21oi_1
XFILLER_31_971 VPWR VGND sg13g2_decap_8
X_4704_ net535 _1527_ mydesign.accum\[60\] _1598_ VPWR VGND sg13g2_nand3_1
XFILLER_33_1015 VPWR VGND sg13g2_decap_8
X_5684_ _2599_ _0384_ net618 _2466_ VPWR VGND sg13g2_nand3_1
X_4635_ net625 VPWR _1538_ VGND net489 _1537_ sg13g2_o21ai_1
X_4566_ _1474_ VPWR _1476_ VGND _1454_ _1456_ sg13g2_o21ai_1
X_3517_ _0543_ _0544_ _0545_ VPWR VGND sg13g2_nor2_1
X_4497_ _1411_ net575 mydesign.pe_weights\[48\] net532 VPWR VGND sg13g2_and3_1
X_3448_ VGND VPWR _0481_ _0489_ _0075_ _0490_ sg13g2_a21oi_1
X_3379_ net622 VPWR _0428_ VGND net1069 net431 sg13g2_o21ai_1
XFILLER_40_1008 VPWR VGND sg13g2_decap_8
X_5118_ _1958_ VPWR _1960_ VGND _1937_ _1939_ sg13g2_o21ai_1
X_6098_ net292 VGND VPWR net750 mydesign.accum\[0\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_5049_ net475 VPWR _1895_ VGND net734 _1894_ sg13g2_o21ai_1
XFILLER_14_949 VPWR VGND sg13g2_decap_8
XFILLER_25_297 VPWR VGND sg13g2_fill_1
X_6028__350 VPWR VGND net350 sg13g2_tiehi
XFILLER_9_419 VPWR VGND sg13g2_fill_1
XFILLER_22_982 VPWR VGND sg13g2_decap_8
XFILLER_49_1000 VPWR VGND sg13g2_decap_8
XFILLER_5_625 VPWR VGND sg13g2_fill_2
XFILLER_49_846 VPWR VGND sg13g2_decap_8
X_5818__124 VPWR VGND net124 sg13g2_tiehi
X_5970__217 VPWR VGND net217 sg13g2_tiehi
XFILLER_48_389 VPWR VGND sg13g2_decap_4
XFILLER_1_1013 VPWR VGND sg13g2_decap_8
XFILLER_16_242 VPWR VGND sg13g2_fill_1
XFILLER_44_562 VPWR VGND sg13g2_decap_8
XFILLER_17_787 VPWR VGND sg13g2_fill_1
XFILLER_16_297 VPWR VGND sg13g2_fill_1
XFILLER_20_919 VPWR VGND sg13g2_decap_8
XFILLER_32_768 VPWR VGND sg13g2_fill_2
X_5825__117 VPWR VGND net117 sg13g2_tiehi
X_4420_ _1346_ mydesign.pe_weights\[54\] mydesign.pe_inputs\[42\] VPWR VGND sg13g2_nand2_1
X_4351_ VGND VPWR _2563_ net440 _0180_ _1288_ sg13g2_a21oi_1
X_6075__112 VPWR VGND net112 sg13g2_tiehi
X_4282_ _1210_ _1224_ _1225_ VPWR VGND sg13g2_and2_1
X_3302_ net788 _2669_ _2691_ _0051_ VPWR VGND sg13g2_mux2_1
X_6021_ net382 VGND VPWR _0247_ mydesign.inputs\[3\]\[7\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_3233_ _2654_ net669 _2650_ VPWR VGND sg13g2_nand2_1
X_3164_ net607 _2597_ _2598_ _2604_ _0000_ VPWR VGND sg13g2_nor4_1
XFILLER_27_507 VPWR VGND sg13g2_fill_2
X_3095_ VPWR _2536_ net943 VGND sg13g2_inv_1
X_3997_ _0968_ VPWR _0972_ VGND _0969_ _0970_ sg13g2_o21ai_1
X_5805_ net143 VGND VPWR _0031_ mydesign.weights\[2\]\[14\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5736_ _2497_ net700 _2495_ VPWR VGND sg13g2_nand2_1
X_5667_ net476 VPWR _2455_ VGND net587 net1049 sg13g2_o21ai_1
X_4618_ mydesign.inputs\[2\]\[17\] mydesign.inputs\[2\]\[13\] net550 _1523_ VPWR VGND
+ sg13g2_mux2_1
X_5598_ _2389_ mydesign.pe_inputs\[5\] mydesign.pe_weights\[18\] VPWR VGND sg13g2_nand2_1
Xhold441 mydesign.accum\[125\] VPWR VGND net1060 sg13g2_dlygate4sd3_1
Xhold463 mydesign.pe_inputs\[46\] VPWR VGND net1082 sg13g2_dlygate4sd3_1
X_4549_ _1459_ mydesign.pe_weights\[49\] mydesign.pe_inputs\[39\] VPWR VGND sg13g2_nand2_1
Xhold430 mydesign.accum\[6\] VPWR VGND net1049 sg13g2_dlygate4sd3_1
Xhold452 mydesign.pe_inputs\[61\] VPWR VGND net1071 sg13g2_dlygate4sd3_1
XFILLER_1_149 VPWR VGND sg13g2_decap_4
Xhold474 mydesign.load_counter\[2\] VPWR VGND net1093 sg13g2_dlygate4sd3_1
Xhold485 _0339_ VPWR VGND net1104 sg13g2_dlygate4sd3_1
XFILLER_46_838 VPWR VGND sg13g2_decap_8
XFILLER_45_337 VPWR VGND sg13g2_decap_4
XFILLER_26_551 VPWR VGND sg13g2_decap_8
XFILLER_14_757 VPWR VGND sg13g2_fill_1
XFILLER_9_216 VPWR VGND sg13g2_decap_4
XFILLER_10_963 VPWR VGND sg13g2_decap_8
XFILLER_49_643 VPWR VGND sg13g2_decap_8
X_3920_ _0906_ _0898_ _0907_ VPWR VGND sg13g2_xor2_1
X_3851_ _0841_ _0838_ _0842_ VPWR VGND sg13g2_xor2_1
XFILLER_32_576 VPWR VGND sg13g2_fill_1
X_3782_ _0779_ VPWR _0780_ VGND net497 mydesign.weights\[2\]\[12\] sg13g2_o21ai_1
X_5521_ _2299_ VPWR _2322_ VGND _2298_ _2301_ sg13g2_o21ai_1
XFILLER_30_1018 VPWR VGND sg13g2_decap_8
X_5452_ net521 mydesign.pe_weights\[20\] net729 _2257_ VPWR VGND _2255_ sg13g2_nand4_1
X_5383_ _2196_ _2188_ _2197_ VPWR VGND sg13g2_xor2_1
X_4403_ _1330_ _1328_ _1329_ VPWR VGND sg13g2_nand2_1
X_4334_ _1256_ _1255_ _1272_ _1274_ VPWR VGND sg13g2_a21o_1
XFILLER_8_1008 VPWR VGND sg13g2_decap_8
X_4265_ VGND VPWR net570 _1207_ _0174_ _1208_ sg13g2_a21oi_1
X_5918__321 VPWR VGND net321 sg13g2_tiehi
X_6004_ net78 VGND VPWR net1032 mydesign.pe_inputs\[26\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_4196_ _1151_ _1152_ _1153_ VPWR VGND sg13g2_nor2b_1
X_3216_ _2643_ VPWR _0013_ VGND net604 _2641_ sg13g2_o21ai_1
X_5863__47 VPWR VGND net47 sg13g2_tiehi
X_3147_ _2588_ net1110 VPWR VGND sg13g2_inv_2
X_3078_ _2519_ net2 VPWR VGND sg13g2_inv_2
X_5719_ _2489_ net614 VPWR VGND _2482_ sg13g2_nand2b_2
Xhold271 mydesign.accum\[29\] VPWR VGND net890 sg13g2_dlygate4sd3_1
Xhold260 mydesign.pe_inputs\[29\] VPWR VGND net879 sg13g2_dlygate4sd3_1
Xhold293 mydesign.accum\[55\] VPWR VGND net912 sg13g2_dlygate4sd3_1
Xhold282 _0238_ VPWR VGND net901 sg13g2_dlygate4sd3_1
XFILLER_49_99 VPWR VGND sg13g2_decap_4
XFILLER_46_635 VPWR VGND sg13g2_decap_8
XFILLER_18_304 VPWR VGND sg13g2_decap_4
X_5815__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_33_307 VPWR VGND sg13g2_decap_8
XFILLER_42_863 VPWR VGND sg13g2_decap_8
XFILLER_14_543 VPWR VGND sg13g2_fill_1
XFILLER_6_764 VPWR VGND sg13g2_fill_1
XFILLER_5_230 VPWR VGND sg13g2_fill_1
XFILLER_2_992 VPWR VGND sg13g2_decap_8
X_4050_ _1001_ _0998_ _1018_ _1022_ VPWR VGND sg13g2_a21o_1
Xinput6 ui_in[6] net6 VPWR VGND sg13g2_buf_2
XFILLER_25_819 VPWR VGND sg13g2_fill_1
X_4952_ _1808_ _1790_ _1807_ VPWR VGND sg13g2_nand2_1
XFILLER_18_882 VPWR VGND sg13g2_fill_2
XFILLER_36_189 VPWR VGND sg13g2_fill_2
X_4883_ _1758_ _1756_ _1757_ VPWR VGND sg13g2_xnor2_1
X_3903_ VGND VPWR net572 _0890_ _0129_ _0891_ sg13g2_a21oi_1
X_3834_ _0826_ _0808_ _0824_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_896 VPWR VGND sg13g2_decap_8
X_5883__383 VPWR VGND net383 sg13g2_tiehi
X_3765_ _0771_ net411 _0770_ VPWR VGND sg13g2_nand2_1
X_5504_ _2305_ VPWR _2306_ VGND _2284_ _2286_ sg13g2_o21ai_1
X_3696_ _0705_ _0706_ _0707_ VPWR VGND sg13g2_nor2b_1
X_5435_ VGND VPWR _2524_ net444 _0308_ _2244_ sg13g2_a21oi_1
XFILLER_0_929 VPWR VGND sg13g2_decap_8
X_5366_ _2181_ _2157_ _2179_ VPWR VGND sg13g2_xnor2_1
X_4317_ _1237_ VPWR _1258_ VGND _1230_ _1238_ sg13g2_o21ai_1
X_5297_ VGND VPWR _2120_ _2121_ _2124_ _2119_ sg13g2_a21oi_1
X_4248_ net471 VPWR _1193_ VGND net570 net983 sg13g2_o21ai_1
X_4179_ _1136_ _1135_ _1137_ VPWR VGND sg13g2_xor2_1
XFILLER_36_690 VPWR VGND sg13g2_fill_1
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
X_6099__284 VPWR VGND net284 sg13g2_tiehi
XFILLER_4_2 VPWR VGND sg13g2_fill_1
XFILLER_3_767 VPWR VGND sg13g2_fill_2
XFILLER_47_922 VPWR VGND sg13g2_decap_8
Xfanout570 net571 net570 VPWR VGND sg13g2_buf_8
Xfanout581 net594 net581 VPWR VGND sg13g2_buf_1
Xfanout592 net593 net592 VPWR VGND sg13g2_buf_8
XFILLER_18_123 VPWR VGND sg13g2_fill_1
XFILLER_20_1017 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_999 VPWR VGND sg13g2_decap_8
XFILLER_14_395 VPWR VGND sg13g2_fill_1
XFILLER_30_899 VPWR VGND sg13g2_decap_8
X_3550_ net468 VPWR _0577_ VGND net559 net1061 sg13g2_o21ai_1
X_5220_ VGND VPWR _2031_ _2047_ _2051_ _2046_ sg13g2_a21oi_1
X_3481_ _0514_ VPWR _0515_ VGND net498 mydesign.weights\[0\]\[20\] sg13g2_o21ai_1
X_5151_ _1991_ _1990_ _1989_ VPWR VGND sg13g2_nand2b_1
X_4102_ VGND VPWR _2576_ net436 _0154_ _1065_ sg13g2_a21oi_1
X_5082_ _1925_ mydesign.pe_weights\[35\] net526 VPWR VGND sg13g2_nand2_1
X_6079__80 VPWR VGND net80 sg13g2_tiehi
X_4033_ VGND VPWR net564 _1005_ _0144_ _1006_ sg13g2_a21oi_1
XFILLER_38_944 VPWR VGND sg13g2_decap_8
X_5984_ net189 VGND VPWR _0210_ mydesign.accum\[70\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_4935_ _1790_ _1791_ _1792_ VPWR VGND sg13g2_nor2b_1
XFILLER_21_811 VPWR VGND sg13g2_decap_4
X_5987__182 VPWR VGND net182 sg13g2_tiehi
X_4866_ _1742_ _1741_ _0241_ VPWR VGND sg13g2_nor2b_1
X_3817_ _0810_ _0808_ _0809_ VPWR VGND sg13g2_nand2_1
X_4797_ _1674_ _1658_ _1677_ VPWR VGND sg13g2_xor2_1
X_3748_ _0756_ _0740_ _0754_ VPWR VGND sg13g2_xnor2_1
X_6022__378 VPWR VGND net378 sg13g2_tiehi
X_3679_ _0690_ mydesign.pe_inputs\[62\] _0648_ VPWR VGND sg13g2_nand2_1
X_5418_ _2212_ _2228_ _2209_ _2230_ VPWR VGND sg13g2_nand3_1
XFILLER_0_715 VPWR VGND sg13g2_decap_4
X_5349_ _2165_ _2149_ _2164_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_944 VPWR VGND sg13g2_decap_8
XFILLER_44_925 VPWR VGND sg13g2_decap_8
XFILLER_46_89 VPWR VGND sg13g2_fill_1
XFILLER_43_413 VPWR VGND sg13g2_decap_8
XFILLER_43_446 VPWR VGND sg13g2_fill_1
XFILLER_12_811 VPWR VGND sg13g2_fill_2
XFILLER_24_671 VPWR VGND sg13g2_fill_2
XFILLER_11_332 VPWR VGND sg13g2_decap_8
XFILLER_11_343 VPWR VGND sg13g2_fill_1
XFILLER_7_39 VPWR VGND sg13g2_fill_2
XFILLER_11_387 VPWR VGND sg13g2_fill_2
XFILLER_4_1011 VPWR VGND sg13g2_decap_8
XFILLER_19_432 VPWR VGND sg13g2_decap_4
XFILLER_46_251 VPWR VGND sg13g2_fill_1
XFILLER_47_796 VPWR VGND sg13g2_decap_8
XFILLER_19_498 VPWR VGND sg13g2_fill_1
XFILLER_35_936 VPWR VGND sg13g2_decap_8
XFILLER_43_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_41_clk clknet_3_4__leaf_clk clknet_leaf_41_clk VPWR VGND sg13g2_buf_8
X_4720_ VGND VPWR _1593_ _1610_ _1613_ _1609_ sg13g2_a21oi_1
X_4651_ _1548_ mydesign.pe_weights\[44\] _1527_ VPWR VGND sg13g2_nand2_1
X_3602_ _0624_ VPWR _0626_ VGND _0610_ _0612_ sg13g2_o21ai_1
X_4582_ _1469_ _1490_ _1491_ VPWR VGND sg13g2_nor2b_1
X_6000__94 VPWR VGND net94 sg13g2_tiehi
X_3533_ net455 _0525_ _2586_ _0560_ VPWR VGND sg13g2_nand3_1
X_3464_ net554 mydesign.inputs\[0\]\[25\] mydesign.inputs\[0\]\[21\] mydesign.inputs\[0\]\[17\]
+ mydesign.inputs\[0\]\[13\] net544 _0501_ VPWR VGND sg13g2_mux4_1
X_5203_ _2035_ mydesign.pe_weights\[28\] _2015_ VPWR VGND sg13g2_nand2_1
X_5134_ _1953_ _1974_ _1975_ VPWR VGND sg13g2_nor2_1
X_3395_ net511 mydesign.accum\[123\] mydesign.accum\[91\] mydesign.accum\[59\] mydesign.accum\[27\]
+ net504 _0442_ VPWR VGND sg13g2_mux4_1
XFILLER_29_207 VPWR VGND sg13g2_fill_2
X_5065_ net526 net530 mydesign.accum\[34\] _1909_ VPWR VGND sg13g2_a21o_1
X_4016_ _0990_ mydesign.pe_inputs\[54\] _0926_ VPWR VGND sg13g2_nand2_1
XFILLER_37_240 VPWR VGND sg13g2_fill_2
XFILLER_16_15 VPWR VGND sg13g2_fill_2
X_5967_ net223 VGND VPWR _0193_ mydesign.accum\[77\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_4918_ VGND VPWR _2537_ net440 _0255_ _1780_ sg13g2_a21oi_1
XFILLER_12_129 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_32_clk clknet_3_5__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
XFILLER_34_991 VPWR VGND sg13g2_decap_8
X_5898_ net357 VGND VPWR net689 mydesign.accum\[104\] clknet_leaf_40_clk sg13g2_dfrbpq_2
XFILLER_21_652 VPWR VGND sg13g2_fill_1
XFILLER_32_14 VPWR VGND sg13g2_fill_2
X_4849_ _1726_ mydesign.pe_weights\[42\] mydesign.pe_inputs\[31\] VPWR VGND sg13g2_nand2_1
XFILLER_10_1005 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_44_722 VPWR VGND sg13g2_decap_8
XFILLER_17_936 VPWR VGND sg13g2_decap_8
XFILLER_28_284 VPWR VGND sg13g2_decap_8
XFILLER_43_221 VPWR VGND sg13g2_fill_2
XFILLER_44_799 VPWR VGND sg13g2_decap_8
XFILLER_43_254 VPWR VGND sg13g2_fill_1
X_6144__200 VPWR VGND net200 sg13g2_tiehi
XFILLER_25_980 VPWR VGND sg13g2_decap_8
XFILLER_43_287 VPWR VGND sg13g2_decap_8
XFILLER_31_449 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_23_clk clknet_3_6__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_40_994 VPWR VGND sg13g2_decap_8
XFILLER_12_685 VPWR VGND sg13g2_fill_1
XFILLER_26_1023 VPWR VGND sg13g2_decap_4
XFILLER_39_516 VPWR VGND sg13g2_fill_2
X_3180_ _2615_ VPWR _0004_ VGND _2608_ _2616_ sg13g2_o21ai_1
XFILLER_35_700 VPWR VGND sg13g2_fill_1
X_5821_ net121 VGND VPWR _0047_ mydesign.inputs\[0\]\[14\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5752_ net612 VPWR _2506_ VGND net985 _2505_ sg13g2_o21ai_1
XFILLER_15_490 VPWR VGND sg13g2_fill_1
XFILLER_16_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_14_clk clknet_3_2__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
XFILLER_31_950 VPWR VGND sg13g2_decap_8
X_4703_ _1597_ mydesign.pe_weights\[46\] _1531_ VPWR VGND sg13g2_nand2b_1
X_5683_ _2465_ VPWR _0335_ VGND net598 _2461_ sg13g2_o21ai_1
X_4634_ _1534_ VPWR _1537_ VGND _1535_ _1536_ sg13g2_o21ai_1
X_4565_ _1454_ _1456_ _1474_ _1475_ VPWR VGND sg13g2_or3_1
X_3516_ _0544_ _0501_ _0520_ VPWR VGND sg13g2_nand2_1
X_4496_ VGND VPWR _2553_ net441 _0203_ _1410_ sg13g2_a21oi_1
X_3447_ net622 VPWR _0490_ VGND net1084 net430 sg13g2_o21ai_1
X_3378_ VPWR VGND net456 _0426_ _0421_ _0405_ _0427_ _0420_ sg13g2_a221oi_1
X_5117_ _1937_ _1939_ _1958_ _1959_ VPWR VGND sg13g2_or3_1
X_6097_ net300 VGND VPWR net681 mydesign.inputs\[3\]\[11\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_5048_ _1894_ net584 mydesign.pe_weights\[32\] net526 VPWR VGND sg13g2_and3_1
XFILLER_14_928 VPWR VGND sg13g2_decap_8
XFILLER_25_265 VPWR VGND sg13g2_fill_2
XFILLER_25_276 VPWR VGND sg13g2_fill_1
XFILLER_40_224 VPWR VGND sg13g2_fill_1
XFILLER_40_213 VPWR VGND sg13g2_decap_8
X_5928__301 VPWR VGND net301 sg13g2_tiehi
XFILLER_40_246 VPWR VGND sg13g2_fill_1
XFILLER_22_961 VPWR VGND sg13g2_decap_8
XFILLER_21_460 VPWR VGND sg13g2_fill_1
XFILLER_5_604 VPWR VGND sg13g2_fill_2
XFILLER_4_158 VPWR VGND sg13g2_fill_2
XFILLER_49_825 VPWR VGND sg13g2_decap_8
XFILLER_1_865 VPWR VGND sg13g2_decap_4
XFILLER_1_887 VPWR VGND sg13g2_decap_8
XFILLER_32_703 VPWR VGND sg13g2_fill_1
XFILLER_40_780 VPWR VGND sg13g2_decap_8
XFILLER_8_420 VPWR VGND sg13g2_fill_1
XFILLER_13_994 VPWR VGND sg13g2_decap_8
XFILLER_9_998 VPWR VGND sg13g2_decap_8
X_4350_ net629 VPWR _1288_ VGND net532 net440 sg13g2_o21ai_1
X_3301_ net766 _2668_ _2691_ _0050_ VPWR VGND sg13g2_mux2_1
XFILLER_4_670 VPWR VGND sg13g2_fill_1
X_4281_ _1223_ _1211_ _1224_ VPWR VGND sg13g2_xor2_1
X_5875__23 VPWR VGND net23 sg13g2_tiehi
X_6020_ net386 VGND VPWR _0246_ mydesign.inputs\[3\]\[6\] clknet_leaf_46_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_3_clk clknet_3_0__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_3232_ _2653_ VPWR _0019_ VGND net600 _2649_ sg13g2_o21ai_1
X_3163_ VPWR _2604_ _2603_ VGND sg13g2_inv_1
X_3094_ VPWR _2535_ net862 VGND sg13g2_inv_1
XFILLER_27_519 VPWR VGND sg13g2_decap_8
X_5804_ net145 VGND VPWR _0030_ mydesign.weights\[2\]\[13\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_35_585 VPWR VGND sg13g2_fill_1
X_3996_ _0968_ _0969_ _0970_ _0971_ VPWR VGND sg13g2_or3_1
X_5735_ _2496_ VPWR _0356_ VGND net604 _2495_ sg13g2_o21ai_1
X_5666_ VGND VPWR _2454_ _2453_ _2452_ sg13g2_or2_1
XFILLER_30_290 VPWR VGND sg13g2_fill_2
XFILLER_31_791 VPWR VGND sg13g2_fill_2
X_4617_ VGND VPWR _2547_ net492 _0212_ _1522_ sg13g2_a21oi_1
X_5597_ _2381_ VPWR _2388_ VGND _2373_ _2382_ sg13g2_o21ai_1
Xhold420 _0314_ VPWR VGND net1039 sg13g2_dlygate4sd3_1
Xhold442 mydesign.accum\[123\] VPWR VGND net1061 sg13g2_dlygate4sd3_1
X_4548_ VGND VPWR net566 _1457_ _0207_ _1458_ sg13g2_a21oi_1
XFILLER_2_607 VPWR VGND sg13g2_fill_1
Xhold453 net14 VPWR VGND net1072 sg13g2_dlygate4sd3_1
Xhold431 mydesign.pe_inputs\[40\] VPWR VGND net1050 sg13g2_dlygate4sd3_1
Xhold464 mydesign.cp\[2\] VPWR VGND net1083 sg13g2_dlygate4sd3_1
X_4479_ VGND VPWR _1401_ _1400_ _2618_ sg13g2_or2_1
Xhold486 mydesign.out\[2\] VPWR VGND net1105 sg13g2_dlygate4sd3_1
Xhold475 mydesign.pe_inputs\[28\] VPWR VGND net1094 sg13g2_dlygate4sd3_1
XFILLER_46_817 VPWR VGND sg13g2_decap_8
X_6149_ net256 VGND VPWR _0375_ mydesign.weights\[1\]\[23\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_22_780 VPWR VGND sg13g2_fill_1
XFILLER_5_412 VPWR VGND sg13g2_decap_8
XFILLER_6_979 VPWR VGND sg13g2_decap_8
XFILLER_5_467 VPWR VGND sg13g2_fill_1
XFILLER_49_622 VPWR VGND sg13g2_decap_8
XFILLER_23_1015 VPWR VGND sg13g2_decap_8
XFILLER_49_699 VPWR VGND sg13g2_decap_8
XFILLER_48_187 VPWR VGND sg13g2_fill_2
XFILLER_17_574 VPWR VGND sg13g2_decap_8
X_3850_ _0839_ mydesign.accum\[107\] _0841_ VPWR VGND sg13g2_xor2_1
X_3781_ VGND VPWR net497 _2589_ _0779_ _0393_ sg13g2_a21oi_1
X_5520_ _2321_ _2316_ _2320_ VPWR VGND sg13g2_xnor2_1
X_5451_ net521 mydesign.pe_weights\[20\] net729 _2256_ VPWR VGND sg13g2_nand3_1
X_4402_ net534 net538 mydesign.accum\[75\] _1329_ VPWR VGND sg13g2_a21o_1
X_5382_ _2196_ _2189_ _2194_ VPWR VGND sg13g2_xnor2_1
X_4333_ _1256_ _1272_ _1255_ _1273_ VPWR VGND sg13g2_nand3_1
X_4264_ net472 VPWR _1208_ VGND net570 net961 sg13g2_o21ai_1
X_3215_ _2643_ net423 _2642_ VPWR VGND sg13g2_nand2_1
X_6003_ net82 VGND VPWR _0229_ mydesign.pe_inputs\[25\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_4195_ VGND VPWR _1152_ _1150_ _1131_ sg13g2_or2_1
XFILLER_39_121 VPWR VGND sg13g2_decap_8
X_6018__394 VPWR VGND net394 sg13g2_tiehi
X_3146_ _2587_ net547 VPWR VGND sg13g2_inv_2
XFILLER_43_809 VPWR VGND sg13g2_decap_8
X_3077_ _2518_ net3 VPWR VGND sg13g2_inv_2
XFILLER_23_500 VPWR VGND sg13g2_fill_2
XFILLER_23_544 VPWR VGND sg13g2_decap_8
XFILLER_23_555 VPWR VGND sg13g2_fill_1
X_3979_ _0953_ _0954_ _0955_ VPWR VGND sg13g2_nor2_1
X_5718_ net777 _2488_ _2481_ _0347_ VPWR VGND sg13g2_mux2_1
X_5649_ _2438_ _2429_ _2437_ VPWR VGND sg13g2_xnor2_1
Xhold261 mydesign.pe_weights\[61\] VPWR VGND net880 sg13g2_dlygate4sd3_1
Xhold250 mydesign.weights\[3\]\[15\] VPWR VGND net869 sg13g2_dlygate4sd3_1
Xhold294 mydesign.accum\[34\] VPWR VGND net913 sg13g2_dlygate4sd3_1
Xhold283 mydesign.accum\[43\] VPWR VGND net902 sg13g2_dlygate4sd3_1
Xhold272 mydesign.pe_weights\[28\] VPWR VGND net891 sg13g2_dlygate4sd3_1
XFILLER_46_614 VPWR VGND sg13g2_decap_8
XFILLER_19_817 VPWR VGND sg13g2_decap_8
XFILLER_19_839 VPWR VGND sg13g2_fill_2
XFILLER_18_327 VPWR VGND sg13g2_fill_2
XFILLER_14_522 VPWR VGND sg13g2_fill_1
XFILLER_26_382 VPWR VGND sg13g2_fill_2
XFILLER_42_842 VPWR VGND sg13g2_decap_8
XFILLER_41_352 VPWR VGND sg13g2_fill_1
XFILLER_14_599 VPWR VGND sg13g2_decap_8
XFILLER_6_710 VPWR VGND sg13g2_fill_1
XFILLER_10_772 VPWR VGND sg13g2_decap_8
XFILLER_6_787 VPWR VGND sg13g2_fill_2
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_2_971 VPWR VGND sg13g2_decap_8
XFILLER_49_485 VPWR VGND sg13g2_decap_8
XFILLER_49_474 VPWR VGND sg13g2_fill_2
XFILLER_37_636 VPWR VGND sg13g2_decap_8
X_4951_ _1807_ _1797_ _1806_ VPWR VGND sg13g2_xnor2_1
X_4882_ _1757_ net912 _1743_ VPWR VGND sg13g2_xnor2_1
X_3902_ net465 VPWR _0891_ VGND net573 net942 sg13g2_o21ai_1
X_3833_ VPWR _0825_ _0824_ VGND sg13g2_inv_1
XFILLER_32_374 VPWR VGND sg13g2_decap_8
X_3764_ net612 _0769_ _0770_ VPWR VGND sg13g2_and2_1
X_5503_ _2304_ _2296_ _2305_ VPWR VGND sg13g2_xor2_1
X_3695_ _0688_ VPWR _0706_ VGND _0702_ _0704_ sg13g2_o21ai_1
X_5434_ net635 VPWR _2244_ VGND net1065 net444 sg13g2_o21ai_1
XFILLER_0_908 VPWR VGND sg13g2_decap_8
X_5365_ _2180_ _2157_ _2179_ VPWR VGND sg13g2_nand2_1
X_4316_ _1256_ _1255_ _1257_ VPWR VGND sg13g2_xor2_1
X_5296_ VGND VPWR net568 _2122_ _0290_ _2123_ sg13g2_a21oi_1
X_4247_ _1190_ _1189_ _1192_ VPWR VGND sg13g2_xor2_1
X_4178_ _1115_ VPWR _1136_ VGND _1096_ _1116_ sg13g2_o21ai_1
X_5844__81 VPWR VGND net81 sg13g2_tiehi
XFILLER_27_102 VPWR VGND sg13g2_fill_1
X_3129_ _2570_ net836 VPWR VGND sg13g2_inv_2
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_23_374 VPWR VGND sg13g2_decap_4
XFILLER_3_702 VPWR VGND sg13g2_decap_8
X_5821__121 VPWR VGND net121 sg13g2_tiehi
Xfanout560 net562 net560 VPWR VGND sg13g2_buf_8
XFILLER_47_901 VPWR VGND sg13g2_decap_8
X_5936__285 VPWR VGND net285 sg13g2_tiehi
Xfanout582 net583 net582 VPWR VGND sg13g2_buf_8
Xfanout571 net595 net571 VPWR VGND sg13g2_buf_8
Xfanout593 net594 net593 VPWR VGND sg13g2_buf_8
XFILLER_18_102 VPWR VGND sg13g2_decap_4
XFILLER_19_647 VPWR VGND sg13g2_decap_4
XFILLER_47_978 VPWR VGND sg13g2_decap_8
XFILLER_46_455 VPWR VGND sg13g2_fill_1
XFILLER_15_831 VPWR VGND sg13g2_fill_1
XFILLER_34_639 VPWR VGND sg13g2_decap_4
XFILLER_14_374 VPWR VGND sg13g2_fill_2
X_3480_ VGND VPWR net498 _2592_ _0514_ net546 sg13g2_a21oi_1
XFILLER_29_1021 VPWR VGND sg13g2_decap_8
X_5150_ _1988_ VPWR _1990_ VGND _1975_ _1978_ sg13g2_o21ai_1
X_4101_ net624 VPWR _1065_ VGND mydesign.pe_weights\[46\] net436 sg13g2_o21ai_1
X_5081_ _1924_ mydesign.pe_weights\[33\] mydesign.pe_inputs\[22\] VPWR VGND sg13g2_nand2_1
XFILLER_38_923 VPWR VGND sg13g2_decap_8
X_4032_ net466 VPWR _1006_ VGND net564 net1006 sg13g2_o21ai_1
XFILLER_49_282 VPWR VGND sg13g2_fill_2
XFILLER_49_271 VPWR VGND sg13g2_fill_2
XFILLER_37_411 VPWR VGND sg13g2_decap_4
X_5983_ net191 VGND VPWR _0209_ mydesign.accum\[69\] clknet_leaf_39_clk sg13g2_dfrbpq_2
XFILLER_25_639 VPWR VGND sg13g2_decap_4
X_4934_ _1789_ VPWR _1791_ VGND _1787_ _1788_ sg13g2_o21ai_1
XFILLER_36_1014 VPWR VGND sg13g2_decap_8
X_4865_ net479 VPWR _1742_ VGND net582 net918 sg13g2_o21ai_1
XFILLER_20_311 VPWR VGND sg13g2_decap_8
XFILLER_21_845 VPWR VGND sg13g2_fill_1
X_3816_ _0789_ mydesign.pe_inputs\[56\] mydesign.accum\[105\] _0809_ VPWR VGND sg13g2_a21o_1
X_4796_ _1658_ _1674_ _1676_ VPWR VGND sg13g2_nor2_1
X_3747_ _0755_ _0754_ _0740_ VPWR VGND sg13g2_nand2b_1
X_3678_ mydesign.pe_inputs\[63\] _0643_ _0689_ VPWR VGND sg13g2_and2_1
X_5417_ VGND VPWR _2209_ _2212_ _2229_ _2228_ sg13g2_a21oi_1
X_5348_ _2164_ _2145_ _2162_ VPWR VGND sg13g2_xnor2_1
X_5279_ _2108_ _2107_ _2106_ VPWR VGND sg13g2_nand2b_1
XFILLER_29_923 VPWR VGND sg13g2_decap_8
XFILLER_44_904 VPWR VGND sg13g2_decap_8
XFILLER_28_466 VPWR VGND sg13g2_fill_2
XFILLER_23_182 VPWR VGND sg13g2_fill_2
XFILLER_8_827 VPWR VGND sg13g2_fill_1
XFILLER_7_315 VPWR VGND sg13g2_decap_8
XFILLER_3_510 VPWR VGND sg13g2_fill_1
XFILLER_11_82 VPWR VGND sg13g2_fill_1
XFILLER_16_8 VPWR VGND sg13g2_decap_8
XFILLER_47_775 VPWR VGND sg13g2_decap_8
XFILLER_35_915 VPWR VGND sg13g2_decap_8
XFILLER_19_477 VPWR VGND sg13g2_fill_1
XFILLER_34_458 VPWR VGND sg13g2_fill_2
XFILLER_36_90 VPWR VGND sg13g2_fill_1
XFILLER_43_970 VPWR VGND sg13g2_decap_8
XFILLER_42_480 VPWR VGND sg13g2_fill_2
XFILLER_30_642 VPWR VGND sg13g2_fill_1
X_4650_ _1547_ _1545_ _1546_ VPWR VGND sg13g2_nand2_1
X_3601_ _0610_ _0612_ _0624_ _0625_ VPWR VGND sg13g2_or3_1
X_4581_ _1488_ _1487_ _1490_ VPWR VGND sg13g2_xor2_1
X_3532_ _0559_ _0501_ _0523_ VPWR VGND sg13g2_nand2_1
X_3463_ net609 _0500_ _0080_ VPWR VGND sg13g2_nor2_1
X_5202_ VGND VPWR net563 _2033_ _0285_ _2034_ sg13g2_a21oi_1
X_5133_ _1974_ _1963_ _1972_ VPWR VGND sg13g2_xnor2_1
X_3394_ VGND VPWR _0405_ _0440_ _0441_ _2698_ sg13g2_a21oi_1
X_5064_ net530 net526 mydesign.accum\[34\] _1908_ VPWR VGND sg13g2_nand3_1
X_4015_ _0989_ _0971_ _0969_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_274 VPWR VGND sg13g2_fill_1
X_5811__131 VPWR VGND net131 sg13g2_tiehi
X_5966_ net225 VGND VPWR _0192_ mydesign.accum\[76\] clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_34_970 VPWR VGND sg13g2_decap_8
X_4917_ net633 VPWR _1780_ VGND mydesign.pe_inputs\[23\] net440 sg13g2_o21ai_1
X_5897_ net359 VGND VPWR _0123_ mydesign.pe_weights\[55\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_4848_ _1712_ VPWR _1725_ VGND _1704_ _1713_ sg13g2_o21ai_1
XFILLER_20_130 VPWR VGND sg13g2_decap_8
X_4779_ _1660_ mydesign.pe_weights\[40\] mydesign.pe_inputs\[29\] VPWR VGND sg13g2_nand2_1
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_535 VPWR VGND sg13g2_fill_2
X_5896__361 VPWR VGND net361 sg13g2_tiehi
XFILLER_48_506 VPWR VGND sg13g2_fill_1
XFILLER_29_720 VPWR VGND sg13g2_fill_2
XFILLER_17_904 VPWR VGND sg13g2_fill_1
XFILLER_29_753 VPWR VGND sg13g2_fill_1
XFILLER_44_701 VPWR VGND sg13g2_decap_8
XFILLER_29_786 VPWR VGND sg13g2_decap_8
XFILLER_29_797 VPWR VGND sg13g2_fill_1
XFILLER_43_211 VPWR VGND sg13g2_decap_4
XFILLER_44_778 VPWR VGND sg13g2_decap_8
XFILLER_32_929 VPWR VGND sg13g2_decap_8
XFILLER_12_631 VPWR VGND sg13g2_fill_1
XFILLER_40_973 VPWR VGND sg13g2_decap_8
XFILLER_12_642 VPWR VGND sg13g2_fill_2
XFILLER_8_646 VPWR VGND sg13g2_fill_2
XFILLER_8_635 VPWR VGND sg13g2_decap_8
XFILLER_12_675 VPWR VGND sg13g2_fill_1
XFILLER_8_657 VPWR VGND sg13g2_fill_2
Xheichips25_template_399 VPWR VGND uio_oe[0] sg13g2_tiehi
X_6040__298 VPWR VGND net298 sg13g2_tiehi
XFILLER_3_362 VPWR VGND sg13g2_fill_2
XFILLER_3_373 VPWR VGND sg13g2_decap_4
XFILLER_26_1002 VPWR VGND sg13g2_decap_8
X_5820_ net122 VGND VPWR _0046_ mydesign.inputs\[0\]\[13\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_16_970 VPWR VGND sg13g2_decap_8
X_5751_ _2591_ _2622_ _2648_ _2505_ VPWR VGND sg13g2_nor3_2
X_4702_ _1578_ VPWR _1596_ VGND _1576_ _1579_ sg13g2_o21ai_1
X_5682_ _2465_ net649 _2461_ VPWR VGND sg13g2_nand2_1
X_4633_ _0392_ VPWR _1536_ VGND net498 mydesign.inputs\[2\]\[15\] sg13g2_o21ai_1
X_4564_ _1472_ _1471_ _1474_ VPWR VGND sg13g2_xor2_1
X_3515_ _0543_ _0541_ _0542_ VPWR VGND sg13g2_nand2_1
X_4495_ net633 VPWR _1410_ VGND net816 net440 sg13g2_o21ai_1
X_3446_ VPWR VGND net456 _0488_ _0483_ net457 _0489_ _0482_ sg13g2_a221oi_1
X_3377_ VGND VPWR net506 _0424_ _0426_ _0425_ sg13g2_a21oi_1
X_5991__146 VPWR VGND net146 sg13g2_tiehi
X_6096_ net308 VGND VPWR net651 mydesign.inputs\[3\]\[10\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_5116_ _1956_ _1955_ _1958_ VPWR VGND sg13g2_xor2_1
X_5047_ VGND VPWR _2529_ net443 _0271_ _1893_ sg13g2_a21oi_1
XFILLER_26_712 VPWR VGND sg13g2_decap_4
XFILLER_26_756 VPWR VGND sg13g2_fill_2
XFILLER_25_255 VPWR VGND sg13g2_fill_2
X_5949_ net259 VGND VPWR _0175_ mydesign.accum\[83\] clknet_leaf_25_clk sg13g2_dfrbpq_2
XFILLER_43_58 VPWR VGND sg13g2_decap_8
XFILLER_22_940 VPWR VGND sg13g2_decap_8
XFILLER_21_483 VPWR VGND sg13g2_fill_1
XFILLER_5_616 VPWR VGND sg13g2_fill_1
XFILLER_0_310 VPWR VGND sg13g2_decap_8
XFILLER_1_822 VPWR VGND sg13g2_decap_8
XFILLER_49_804 VPWR VGND sg13g2_decap_8
XFILLER_0_354 VPWR VGND sg13g2_decap_8
XFILLER_0_376 VPWR VGND sg13g2_decap_8
XFILLER_17_712 VPWR VGND sg13g2_fill_1
XFILLER_16_266 VPWR VGND sg13g2_fill_2
XFILLER_32_737 VPWR VGND sg13g2_decap_4
XFILLER_8_410 VPWR VGND sg13g2_fill_1
XFILLER_9_933 VPWR VGND sg13g2_fill_2
XFILLER_12_450 VPWR VGND sg13g2_fill_1
XFILLER_13_973 VPWR VGND sg13g2_decap_8
XFILLER_9_977 VPWR VGND sg13g2_decap_8
XFILLER_4_660 VPWR VGND sg13g2_fill_1
X_3300_ net780 _2667_ _2691_ _0049_ VPWR VGND sg13g2_mux2_1
X_4280_ _1223_ _1199_ _1221_ VPWR VGND sg13g2_xnor2_1
X_3231_ _2653_ net704 _2650_ VPWR VGND sg13g2_nand2_1
X_3162_ net499 _2600_ _2603_ VPWR VGND sg13g2_nor2_2
XFILLER_48_881 VPWR VGND sg13g2_decap_8
X_3093_ VPWR _2534_ net830 VGND sg13g2_inv_1
XFILLER_23_704 VPWR VGND sg13g2_fill_2
X_5803_ net147 VGND VPWR _0029_ mydesign.weights\[2\]\[12\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_23_726 VPWR VGND sg13g2_fill_1
X_3995_ VGND VPWR mydesign.pe_inputs\[52\] net428 _0970_ mydesign.accum\[99\] sg13g2_a21oi_1
XFILLER_23_759 VPWR VGND sg13g2_decap_4
X_5734_ _2496_ net647 _2495_ VPWR VGND sg13g2_nand2_1
X_5665_ VGND VPWR _2439_ _2441_ _2453_ _2451_ sg13g2_a21oi_1
X_4616_ net624 VPWR _1522_ VGND net485 _1521_ sg13g2_o21ai_1
X_5596_ _2387_ net1111 mydesign.pe_weights\[19\] VPWR VGND sg13g2_nand2_1
Xhold410 mydesign.accum\[17\] VPWR VGND net1029 sg13g2_dlygate4sd3_1
Xhold443 mydesign.accum\[126\] VPWR VGND net1062 sg13g2_dlygate4sd3_1
Xhold421 mydesign.accum\[2\] VPWR VGND net1040 sg13g2_dlygate4sd3_1
X_4547_ net464 VPWR _1458_ VGND net566 net906 sg13g2_o21ai_1
Xhold454 mydesign.pe_inputs\[56\] VPWR VGND net1073 sg13g2_dlygate4sd3_1
Xhold432 _0164_ VPWR VGND net1051 sg13g2_dlygate4sd3_1
Xhold476 mydesign.pe_inputs\[36\] VPWR VGND net1095 sg13g2_dlygate4sd3_1
Xhold487 mydesign.load_counter\[1\] VPWR VGND net1106 sg13g2_dlygate4sd3_1
X_4478_ _1400_ _2619_ _2607_ VPWR VGND sg13g2_nand2b_1
Xhold465 net15 VPWR VGND net1084 sg13g2_dlygate4sd3_1
X_3429_ mydesign.accum\[118\] mydesign.accum\[86\] net512 _0473_ VPWR VGND sg13g2_mux2_1
X_6148_ net272 VGND VPWR _0374_ mydesign.weights\[1\]\[22\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_6079_ net80 VGND VPWR _0305_ mydesign.accum\[21\] clknet_leaf_26_clk sg13g2_dfrbpq_2
XFILLER_26_520 VPWR VGND sg13g2_decap_4
XFILLER_26_586 VPWR VGND sg13g2_fill_2
XFILLER_16_1012 VPWR VGND sg13g2_decap_8
X_6141__248 VPWR VGND net248 sg13g2_tiehi
XFILLER_22_792 VPWR VGND sg13g2_fill_2
XFILLER_6_936 VPWR VGND sg13g2_decap_4
XFILLER_5_402 VPWR VGND sg13g2_decap_4
XFILLER_6_958 VPWR VGND sg13g2_decap_8
XFILLER_10_998 VPWR VGND sg13g2_decap_8
X_5902__349 VPWR VGND net349 sg13g2_tiehi
XFILLER_49_601 VPWR VGND sg13g2_decap_8
XFILLER_49_678 VPWR VGND sg13g2_decap_8
XFILLER_45_884 VPWR VGND sg13g2_decap_8
XFILLER_32_556 VPWR VGND sg13g2_fill_2
XFILLER_32_567 VPWR VGND sg13g2_decap_8
X_3780_ VGND VPWR _2580_ net435 _0119_ _0778_ sg13g2_a21oi_1
X_5946__265 VPWR VGND net265 sg13g2_tiehi
X_5450_ _2253_ _2254_ _2255_ VPWR VGND sg13g2_nor2b_1
X_4401_ net538 mydesign.pe_inputs\[40\] mydesign.accum\[75\] _1328_ VPWR VGND sg13g2_nand3_1
X_5381_ _2195_ _2189_ _2194_ VPWR VGND sg13g2_nand2_1
X_4332_ _1272_ _1269_ _1270_ VPWR VGND sg13g2_xnor2_1
X_5799__151 VPWR VGND net151 sg13g2_tiehi
X_4263_ _1207_ _1191_ _1206_ VPWR VGND sg13g2_xnor2_1
X_3214_ VGND VPWR net609 _2642_ _2640_ net605 sg13g2_a21oi_2
X_6002_ net86 VGND VPWR net1023 mydesign.pe_inputs\[24\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_4194_ _1131_ _1150_ _1151_ VPWR VGND sg13g2_and2_1
XFILLER_39_166 VPWR VGND sg13g2_fill_1
XFILLER_39_155 VPWR VGND sg13g2_decap_8
X_3145_ net541 _2586_ VPWR VGND sg13g2_inv_4
X_3076_ _2517_ net4 VPWR VGND sg13g2_inv_2
XFILLER_39_1012 VPWR VGND sg13g2_decap_8
XFILLER_23_512 VPWR VGND sg13g2_fill_1
XFILLER_35_361 VPWR VGND sg13g2_fill_2
XFILLER_36_895 VPWR VGND sg13g2_decap_8
X_3978_ _0954_ _0950_ _0952_ _0919_ mydesign.pe_inputs\[53\] VPWR VGND sg13g2_a22oi_1
X_5717_ _2517_ _2484_ _2488_ VPWR VGND sg13g2_nor2_2
X_5648_ _2434_ _2430_ _2437_ VPWR VGND sg13g2_xor2_1
X_5579_ net475 VPWR _2372_ VGND net587 net1057 sg13g2_o21ai_1
Xhold262 mydesign.pe_weights\[63\] VPWR VGND net881 sg13g2_dlygate4sd3_1
Xhold240 _1772_ VPWR VGND net859 sg13g2_dlygate4sd3_1
XFILLER_2_416 VPWR VGND sg13g2_fill_2
Xhold251 _2509_ VPWR VGND net870 sg13g2_dlygate4sd3_1
XFILLER_49_35 VPWR VGND sg13g2_decap_4
XFILLER_46_1027 VPWR VGND sg13g2_fill_2
Xhold295 _0274_ VPWR VGND net914 sg13g2_dlygate4sd3_1
Xhold284 mydesign.pe_weights\[16\] VPWR VGND net903 sg13g2_dlygate4sd3_1
Xhold273 mydesign.accum\[49\] VPWR VGND net892 sg13g2_dlygate4sd3_1
XFILLER_14_501 VPWR VGND sg13g2_decap_4
XFILLER_26_350 VPWR VGND sg13g2_decap_4
XFILLER_26_394 VPWR VGND sg13g2_decap_8
XFILLER_42_898 VPWR VGND sg13g2_decap_8
XFILLER_5_298 VPWR VGND sg13g2_decap_8
XFILLER_2_950 VPWR VGND sg13g2_decap_8
XFILLER_39_7 VPWR VGND sg13g2_fill_2
XFILLER_36_125 VPWR VGND sg13g2_fill_2
XFILLER_45_681 VPWR VGND sg13g2_decap_8
X_4950_ _1803_ _1787_ _1806_ VPWR VGND sg13g2_xor2_1
XFILLER_18_884 VPWR VGND sg13g2_fill_1
X_4881_ VGND VPWR _1732_ _1747_ _1756_ _1746_ sg13g2_a21oi_1
X_3901_ _0890_ _0876_ _0889_ VPWR VGND sg13g2_xnor2_1
X_3832_ _0824_ _0821_ _0822_ VPWR VGND sg13g2_xnor2_1
X_3763_ _2638_ _2647_ net610 _0769_ VPWR VGND sg13g2_nand3_1
X_5502_ _2304_ _2297_ _2302_ VPWR VGND sg13g2_xnor2_1
X_3694_ _0688_ _0702_ _0704_ _0705_ VPWR VGND sg13g2_nor3_1
X_5433_ VGND VPWR net593 _2242_ _0307_ _2243_ sg13g2_a21oi_1
X_5364_ _2177_ _2170_ _2179_ VPWR VGND sg13g2_xor2_1
X_4315_ _1233_ VPWR _1256_ VGND _1232_ _1235_ sg13g2_o21ai_1
X_5295_ net470 VPWR _2123_ VGND net568 net945 sg13g2_o21ai_1
X_4246_ mydesign.pe_weights\[56\] net536 net739 _1191_ VPWR VGND _1189_ sg13g2_nand4_1
X_4177_ _1135_ _1134_ _1133_ VPWR VGND sg13g2_nand2b_1
X_3128_ VPWR _2569_ net1082 VGND sg13g2_inv_1
XFILLER_27_136 VPWR VGND sg13g2_decap_8
XFILLER_27_147 VPWR VGND sg13g2_fill_1
XFILLER_24_876 VPWR VGND sg13g2_decap_8
X_6013__38 VPWR VGND net38 sg13g2_tiehi
XFILLER_11_526 VPWR VGND sg13g2_decap_8
XFILLER_13_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_725 VPWR VGND sg13g2_fill_2
XFILLER_3_769 VPWR VGND sg13g2_fill_1
XFILLER_3_758 VPWR VGND sg13g2_decap_4
Xfanout550 net552 net550 VPWR VGND sg13g2_buf_8
Xfanout561 net562 net561 VPWR VGND sg13g2_buf_1
Xfanout572 net573 net572 VPWR VGND sg13g2_buf_8
Xfanout583 net594 net583 VPWR VGND sg13g2_buf_8
XFILLER_47_957 VPWR VGND sg13g2_decap_8
Xfanout594 net595 net594 VPWR VGND sg13g2_buf_8
XFILLER_33_139 VPWR VGND sg13g2_fill_2
X_5789__161 VPWR VGND net161 sg13g2_tiehi
XFILLER_25_70 VPWR VGND sg13g2_decap_8
XFILLER_41_183 VPWR VGND sg13g2_fill_2
XFILLER_29_1000 VPWR VGND sg13g2_decap_8
X_4100_ VGND VPWR _2577_ net436 _0153_ _1064_ sg13g2_a21oi_1
X_5080_ _1923_ mydesign.pe_weights\[32\] mydesign.pe_inputs\[23\] VPWR VGND sg13g2_nand2_1
X_5796__154 VPWR VGND net154 sg13g2_tiehi
XFILLER_38_902 VPWR VGND sg13g2_decap_8
X_4031_ _1003_ _1002_ _1005_ VPWR VGND sg13g2_xor2_1
XFILLER_38_979 VPWR VGND sg13g2_decap_8
X_5982_ net193 VGND VPWR _0208_ mydesign.accum\[68\] clknet_leaf_39_clk sg13g2_dfrbpq_2
XFILLER_18_670 VPWR VGND sg13g2_fill_1
X_4933_ _1787_ _1788_ _1789_ _1790_ VPWR VGND sg13g2_nor3_1
XFILLER_18_692 VPWR VGND sg13g2_fill_2
XFILLER_24_139 VPWR VGND sg13g2_fill_2
X_4864_ net582 VPWR _1741_ VGND _1739_ _1740_ sg13g2_o21ai_1
XFILLER_33_684 VPWR VGND sg13g2_fill_2
XFILLER_33_695 VPWR VGND sg13g2_fill_2
X_3815_ mydesign.pe_inputs\[56\] _0789_ mydesign.accum\[105\] _0808_ VPWR VGND sg13g2_nand3_1
X_4795_ _1675_ _1658_ _1674_ VPWR VGND sg13g2_nand2_1
X_3746_ _0754_ _0738_ _0752_ VPWR VGND sg13g2_xnor2_1
X_6003__82 VPWR VGND net82 sg13g2_tiehi
X_5416_ _2228_ _2226_ _2227_ VPWR VGND sg13g2_nand2_1
X_3677_ VGND VPWR _0664_ _0679_ _0688_ _0681_ sg13g2_a21oi_1
X_5347_ _2163_ _2145_ _2162_ VPWR VGND sg13g2_nand2_1
XFILLER_43_1019 VPWR VGND sg13g2_decap_8
XFILLER_0_739 VPWR VGND sg13g2_decap_4
X_5278_ VGND VPWR _2107_ _2105_ _2088_ sg13g2_or2_1
X_4229_ VGND VPWR _2567_ net447 _0168_ _1178_ sg13g2_a21oi_1
XFILLER_46_14 VPWR VGND sg13g2_fill_1
XFILLER_29_979 VPWR VGND sg13g2_decap_8
XFILLER_28_489 VPWR VGND sg13g2_decap_8
XFILLER_12_813 VPWR VGND sg13g2_fill_1
XFILLER_24_673 VPWR VGND sg13g2_fill_1
XFILLER_7_305 VPWR VGND sg13g2_fill_1
XFILLER_7_327 VPWR VGND sg13g2_decap_8
XFILLER_20_890 VPWR VGND sg13g2_fill_1
XFILLER_11_72 VPWR VGND sg13g2_fill_1
XFILLER_47_754 VPWR VGND sg13g2_decap_8
XFILLER_46_242 VPWR VGND sg13g2_decap_8
XFILLER_34_426 VPWR VGND sg13g2_fill_1
XFILLER_14_161 VPWR VGND sg13g2_fill_1
X_3600_ _0624_ _0608_ _0622_ VPWR VGND sg13g2_xnor2_1
X_4580_ _1489_ _1487_ _1488_ VPWR VGND sg13g2_nand2_1
X_3531_ _0558_ _0506_ _0520_ VPWR VGND sg13g2_nand2_1
XFILLER_7_894 VPWR VGND sg13g2_decap_8
X_3462_ _0500_ net455 _0499_ net484 net540 VPWR VGND sg13g2_a22oi_1
X_5201_ net466 VPWR _2034_ VGND net563 net954 sg13g2_o21ai_1
X_3393_ net515 mydesign.accum\[115\] mydesign.accum\[83\] mydesign.accum\[51\] mydesign.accum\[19\]
+ net508 _0440_ VPWR VGND sg13g2_mux4_1
X_5132_ _1973_ _1963_ _1972_ VPWR VGND sg13g2_nand2_1
XFILLER_28_0 VPWR VGND sg13g2_fill_2
X_5063_ _1907_ mydesign.pe_weights\[33\] mydesign.pe_inputs\[21\] VPWR VGND sg13g2_nand2_1
XFILLER_38_765 VPWR VGND sg13g2_decap_8
X_4014_ _0988_ mydesign.pe_inputs\[55\] _0919_ VPWR VGND sg13g2_nand2_1
XFILLER_16_17 VPWR VGND sg13g2_fill_1
XFILLER_25_404 VPWR VGND sg13g2_decap_8
XFILLER_25_415 VPWR VGND sg13g2_fill_1
XFILLER_19_990 VPWR VGND sg13g2_decap_8
X_5965_ net227 VGND VPWR _0191_ mydesign.accum\[75\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_4916_ VGND VPWR _2538_ net442 _0254_ _1779_ sg13g2_a21oi_1
X_5896_ net361 VGND VPWR _0122_ mydesign.pe_weights\[54\] clknet_leaf_41_clk sg13g2_dfrbpq_2
X_4847_ _1723_ _1724_ _0240_ VPWR VGND sg13g2_nor2_1
X_4778_ VGND VPWR mydesign.pe_weights\[41\] net529 _1659_ mydesign.accum\[49\] sg13g2_a21oi_1
X_3729_ _0738_ _0736_ _0737_ VPWR VGND sg13g2_nand2b_1
XFILLER_0_514 VPWR VGND sg13g2_decap_8
XFILLER_28_231 VPWR VGND sg13g2_fill_1
XFILLER_44_757 VPWR VGND sg13g2_decap_8
XFILLER_43_223 VPWR VGND sg13g2_fill_1
XFILLER_16_459 VPWR VGND sg13g2_decap_4
XFILLER_32_908 VPWR VGND sg13g2_decap_8
XFILLER_40_952 VPWR VGND sg13g2_decap_8
X_5793__157 VPWR VGND net157 sg13g2_tiehi
XFILLER_47_551 VPWR VGND sg13g2_decap_8
XFILLER_19_264 VPWR VGND sg13g2_fill_2
XFILLER_34_223 VPWR VGND sg13g2_decap_8
X_5750_ _2504_ VPWR _0363_ VGND _1775_ _2500_ sg13g2_o21ai_1
XFILLER_30_440 VPWR VGND sg13g2_fill_1
X_5681_ _2464_ VPWR _0334_ VGND net600 _2461_ sg13g2_o21ai_1
X_4701_ _1595_ mydesign.pe_weights\[45\] _1537_ VPWR VGND sg13g2_nand2_1
X_4632_ net557 mydesign.inputs\[2\]\[19\] _1535_ VPWR VGND sg13g2_nor2_1
XFILLER_31_985 VPWR VGND sg13g2_decap_8
X_4563_ _1473_ _1471_ _1472_ VPWR VGND sg13g2_nand2_1
XFILLER_7_680 VPWR VGND sg13g2_fill_1
X_4494_ VGND VPWR _2554_ net440 _0202_ _1409_ sg13g2_a21oi_1
X_3514_ _0523_ _0498_ mydesign.accum\[122\] _0542_ VPWR VGND sg13g2_a21o_1
X_3445_ VGND VPWR net509 _0486_ _0488_ _0487_ sg13g2_a21oi_1
X_5956__245 VPWR VGND net245 sg13g2_tiehi
X_3376_ _0412_ VPWR _0425_ VGND net507 _0422_ sg13g2_o21ai_1
X_5115_ _1957_ _1955_ _1956_ VPWR VGND sg13g2_nand2_1
X_6095_ net316 VGND VPWR net659 mydesign.inputs\[3\]\[9\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_5046_ net634 VPWR _1893_ VGND mydesign.pe_weights\[19\] net442 sg13g2_o21ai_1
XFILLER_26_724 VPWR VGND sg13g2_fill_2
XFILLER_41_727 VPWR VGND sg13g2_fill_1
X_5948_ net261 VGND VPWR net962 mydesign.accum\[82\] clknet_leaf_25_clk sg13g2_dfrbpq_2
XFILLER_22_996 VPWR VGND sg13g2_decap_8
X_5879_ net391 VGND VPWR net852 mydesign.accum\[113\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_5_606 VPWR VGND sg13g2_fill_1
XFILLER_49_1014 VPWR VGND sg13g2_decap_8
XFILLER_1_801 VPWR VGND sg13g2_decap_8
XFILLER_48_304 VPWR VGND sg13g2_fill_1
XFILLER_1_1027 VPWR VGND sg13g2_fill_2
XFILLER_44_543 VPWR VGND sg13g2_fill_2
XFILLER_16_278 VPWR VGND sg13g2_fill_2
XFILLER_16_289 VPWR VGND sg13g2_fill_1
XFILLER_17_93 VPWR VGND sg13g2_decap_8
XFILLER_13_952 VPWR VGND sg13g2_decap_8
XFILLER_12_473 VPWR VGND sg13g2_fill_1
X_3230_ _2652_ VPWR _0018_ VGND net602 _2649_ sg13g2_o21ai_1
X_3161_ _2602_ net563 _2591_ VPWR VGND sg13g2_nand2_2
XFILLER_48_860 VPWR VGND sg13g2_decap_8
X_3092_ VPWR _2533_ net531 VGND sg13g2_inv_1
XFILLER_35_521 VPWR VGND sg13g2_fill_1
XFILLER_35_554 VPWR VGND sg13g2_decap_8
X_5802_ net148 VGND VPWR _0028_ mydesign.inputs\[1\]\[15\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_35_576 VPWR VGND sg13g2_decap_4
X_3994_ _0969_ mydesign.accum\[99\] mydesign.pe_inputs\[52\] net428 VPWR VGND sg13g2_and3_1
XFILLER_22_237 VPWR VGND sg13g2_decap_8
X_5733_ _2495_ net462 _2686_ VPWR VGND sg13g2_nand2_2
X_5664_ _2452_ _2439_ _2441_ _2451_ VPWR VGND sg13g2_and3_1
X_5595_ VGND VPWR net586 _2385_ _0326_ _2386_ sg13g2_a21oi_1
X_4615_ VGND VPWR _1521_ _1520_ _1517_ sg13g2_or2_1
X_4546_ _1455_ _1438_ _1457_ VPWR VGND sg13g2_xor2_1
Xhold400 mydesign.accum\[45\] VPWR VGND net1019 sg13g2_dlygate4sd3_1
Xhold411 _0301_ VPWR VGND net1030 sg13g2_dlygate4sd3_1
Xhold422 _0326_ VPWR VGND net1041 sg13g2_dlygate4sd3_1
Xhold444 mydesign.accum\[5\] VPWR VGND net1063 sg13g2_dlygate4sd3_1
Xhold433 mydesign.accum\[14\] VPWR VGND net1052 sg13g2_dlygate4sd3_1
Xhold477 mydesign.pe_weights\[59\] VPWR VGND net1096 sg13g2_dlygate4sd3_1
Xhold455 _0096_ VPWR VGND net1074 sg13g2_dlygate4sd3_1
Xhold466 _0075_ VPWR VGND net1085 sg13g2_dlygate4sd3_1
X_4477_ VGND VPWR net581 _1398_ _0195_ _1399_ sg13g2_a21oi_1
X_3428_ net513 mydesign.accum\[102\] mydesign.accum\[70\] mydesign.accum\[38\] mydesign.accum\[6\]
+ net506 _0472_ VPWR VGND sg13g2_mux4_1
Xhold488 mydesign.pe_inputs\[20\] VPWR VGND net1107 sg13g2_dlygate4sd3_1
X_3359_ mydesign.accum\[104\] mydesign.accum\[72\] net514 _0409_ VPWR VGND sg13g2_mux2_1
X_6147_ net288 VGND VPWR _0373_ mydesign.weights\[1\]\[21\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_6078_ net88 VGND VPWR _0304_ mydesign.accum\[20\] clknet_leaf_27_clk sg13g2_dfrbpq_2
XFILLER_39_893 VPWR VGND sg13g2_decap_8
XFILLER_38_370 VPWR VGND sg13g2_fill_2
X_5029_ _1879_ VPWR _1881_ VGND _1865_ _1868_ sg13g2_o21ai_1
XFILLER_26_565 VPWR VGND sg13g2_fill_1
XFILLER_14_738 VPWR VGND sg13g2_fill_2
XFILLER_14_749 VPWR VGND sg13g2_fill_1
XFILLER_22_760 VPWR VGND sg13g2_fill_1
XFILLER_10_933 VPWR VGND sg13g2_decap_8
XFILLER_10_977 VPWR VGND sg13g2_decap_8
XFILLER_49_657 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_fill_1
XFILLER_45_863 VPWR VGND sg13g2_decap_8
XFILLER_13_760 VPWR VGND sg13g2_fill_2
XFILLER_8_230 VPWR VGND sg13g2_decap_4
X_4400_ _1327_ mydesign.pe_weights\[54\] mydesign.pe_inputs\[41\] VPWR VGND sg13g2_nand2_1
X_5380_ _2193_ _2190_ _2194_ VPWR VGND sg13g2_xor2_1
X_4331_ VPWR _1271_ _1270_ VGND sg13g2_inv_1
X_4262_ _1206_ _1187_ _1204_ VPWR VGND sg13g2_xnor2_1
X_6001_ net90 VGND VPWR _0227_ mydesign.accum\[63\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3213_ _2641_ net606 _2640_ VPWR VGND sg13g2_nand2_2
X_4193_ _1150_ _1140_ _1148_ VPWR VGND sg13g2_xnor2_1
X_3144_ VPWR _2585_ net756 VGND sg13g2_inv_1
X_3075_ net590 _2516_ VPWR VGND sg13g2_inv_4
XFILLER_36_863 VPWR VGND sg13g2_decap_4
XFILLER_35_351 VPWR VGND sg13g2_fill_2
XFILLER_35_395 VPWR VGND sg13g2_decap_8
X_3977_ mydesign.pe_inputs\[53\] _0919_ _0950_ _0952_ _0953_ VPWR VGND sg13g2_and4_1
X_5716_ net770 _2487_ _2481_ _0346_ VPWR VGND sg13g2_mux2_1
X_5808__137 VPWR VGND net137 sg13g2_tiehi
X_5647_ _2430_ _2434_ _2436_ VPWR VGND sg13g2_nor2_1
XFILLER_3_907 VPWR VGND sg13g2_fill_1
X_5578_ _2369_ _2368_ _2371_ VPWR VGND sg13g2_xor2_1
XFILLER_46_1006 VPWR VGND sg13g2_decap_8
X_4529_ _1440_ mydesign.pe_weights\[48\] mydesign.pe_inputs\[39\] VPWR VGND sg13g2_nand2_1
Xhold241 _0249_ VPWR VGND net860 sg13g2_dlygate4sd3_1
Xhold252 _0367_ VPWR VGND net871 sg13g2_dlygate4sd3_1
Xhold230 mydesign.pe_inputs\[25\] VPWR VGND net849 sg13g2_dlygate4sd3_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
Xhold296 mydesign.accum\[22\] VPWR VGND net915 sg13g2_dlygate4sd3_1
Xhold285 _0268_ VPWR VGND net904 sg13g2_dlygate4sd3_1
Xhold263 mydesign.accum\[74\] VPWR VGND net882 sg13g2_dlygate4sd3_1
Xhold274 _0237_ VPWR VGND net893 sg13g2_dlygate4sd3_1
XFILLER_49_69 VPWR VGND sg13g2_decap_8
XFILLER_46_649 VPWR VGND sg13g2_decap_8
XFILLER_42_877 VPWR VGND sg13g2_decap_8
XFILLER_14_579 VPWR VGND sg13g2_decap_4
XFILLER_2_940 VPWR VGND sg13g2_fill_1
XFILLER_49_465 VPWR VGND sg13g2_fill_1
XFILLER_49_454 VPWR VGND sg13g2_decap_8
X_5999__98 VPWR VGND net98 sg13g2_tiehi
XFILLER_36_137 VPWR VGND sg13g2_decap_4
XFILLER_45_660 VPWR VGND sg13g2_decap_8
X_4880_ _1752_ VPWR _1755_ VGND _1735_ _1748_ sg13g2_o21ai_1
X_3900_ _0889_ _0868_ _0887_ VPWR VGND sg13g2_xnor2_1
X_3831_ _0823_ mydesign.pe_inputs\[57\] _0789_ _0821_ VPWR VGND sg13g2_and3_2
X_3762_ VGND VPWR net570 _0767_ _0111_ _0768_ sg13g2_a21oi_1
XFILLER_20_549 VPWR VGND sg13g2_fill_1
XFILLER_9_561 VPWR VGND sg13g2_fill_1
X_5501_ _2303_ _2297_ _2302_ VPWR VGND sg13g2_nand2_1
X_3693_ VGND VPWR _0700_ _0701_ _0704_ _0689_ sg13g2_a21oi_1
X_5432_ net482 VPWR _2243_ VGND net593 net978 sg13g2_o21ai_1
X_5363_ _2170_ _2177_ _2178_ VPWR VGND sg13g2_nor2_1
X_4314_ _1255_ _1250_ _1254_ VPWR VGND sg13g2_xnor2_1
X_5294_ _2122_ _2120_ _2121_ VPWR VGND sg13g2_xnor2_1
X_4245_ mydesign.pe_weights\[56\] net536 net739 _1190_ VPWR VGND sg13g2_nand3_1
X_4176_ _1112_ _1132_ _1110_ _1134_ VPWR VGND sg13g2_nand3_1
X_3127_ _2568_ net956 VPWR VGND sg13g2_inv_2
XFILLER_28_638 VPWR VGND sg13g2_decap_4
Xfanout551 net552 net551 VPWR VGND sg13g2_buf_1
Xfanout540 net1102 net540 VPWR VGND sg13g2_buf_8
Xfanout562 net595 net562 VPWR VGND sg13g2_buf_2
Xfanout584 net585 net584 VPWR VGND sg13g2_buf_8
Xfanout573 net576 net573 VPWR VGND sg13g2_buf_8
XFILLER_47_936 VPWR VGND sg13g2_decap_8
XFILLER_46_413 VPWR VGND sg13g2_decap_8
Xfanout595 net867 net595 VPWR VGND sg13g2_buf_8
XFILLER_19_638 VPWR VGND sg13g2_fill_2
XFILLER_18_137 VPWR VGND sg13g2_fill_1
X_6147__288 VPWR VGND net288 sg13g2_tiehi
X_6043__286 VPWR VGND net286 sg13g2_tiehi
X_4030_ _1004_ _1002_ _1003_ VPWR VGND sg13g2_nand2b_1
XFILLER_1_280 VPWR VGND sg13g2_fill_2
X_5915__327 VPWR VGND net327 sg13g2_tiehi
XFILLER_38_958 VPWR VGND sg13g2_decap_8
XFILLER_37_446 VPWR VGND sg13g2_decap_4
XFILLER_37_468 VPWR VGND sg13g2_decap_4
X_5981_ net195 VGND VPWR _0207_ mydesign.accum\[67\] clknet_leaf_45_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_44_clk clknet_3_4__leaf_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
X_4932_ _1789_ mydesign.pe_weights\[36\] mydesign.pe_inputs\[25\] VPWR VGND sg13g2_nand2_1
XFILLER_17_192 VPWR VGND sg13g2_fill_2
XFILLER_33_641 VPWR VGND sg13g2_fill_2
X_4863_ VGND VPWR _1719_ _1722_ _1740_ _1738_ sg13g2_a21oi_1
XFILLER_20_324 VPWR VGND sg13g2_decap_8
X_3814_ VGND VPWR net688 _0806_ _0124_ _0807_ sg13g2_a21oi_1
XFILLER_32_195 VPWR VGND sg13g2_decap_8
X_4794_ _1672_ _1669_ _1674_ VPWR VGND sg13g2_xor2_1
X_3745_ _0753_ _0752_ _0738_ VPWR VGND sg13g2_nand2b_1
X_5415_ mydesign.pe_weights\[27\] mydesign.pe_inputs\[15\] mydesign.accum\[22\] _2227_
+ VPWR VGND sg13g2_a21o_1
X_3676_ _0683_ VPWR _0687_ VGND _0669_ _0684_ sg13g2_o21ai_1
X_5994__134 VPWR VGND net134 sg13g2_tiehi
X_5346_ _2162_ _2152_ _2161_ VPWR VGND sg13g2_xnor2_1
X_5277_ _2088_ _2105_ _2106_ VPWR VGND sg13g2_and2_1
XFILLER_29_903 VPWR VGND sg13g2_fill_2
X_4228_ net631 VPWR _1178_ VGND net1013 net447 sg13g2_o21ai_1
X_4159_ _1118_ _1096_ _1117_ VPWR VGND sg13g2_xnor2_1
XFILLER_46_59 VPWR VGND sg13g2_fill_1
XFILLER_29_958 VPWR VGND sg13g2_decap_8
XFILLER_44_939 VPWR VGND sg13g2_decap_8
XFILLER_37_980 VPWR VGND sg13g2_decap_8
XFILLER_15_107 VPWR VGND sg13g2_decap_4
XFILLER_28_468 VPWR VGND sg13g2_fill_1
XFILLER_15_129 VPWR VGND sg13g2_fill_2
XFILLER_36_490 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_35_clk clknet_3_5__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_12_803 VPWR VGND sg13g2_fill_2
X_5966__225 VPWR VGND net225 sg13g2_tiehi
XFILLER_8_818 VPWR VGND sg13g2_decap_8
XFILLER_11_357 VPWR VGND sg13g2_fill_2
XFILLER_11_368 VPWR VGND sg13g2_decap_8
XFILLER_3_545 VPWR VGND sg13g2_fill_1
XFILLER_3_556 VPWR VGND sg13g2_fill_1
XFILLER_4_1025 VPWR VGND sg13g2_decap_4
XFILLER_47_733 VPWR VGND sg13g2_decap_8
XFILLER_28_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_26_clk clknet_3_7__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_30_677 VPWR VGND sg13g2_fill_2
X_3530_ _0557_ _0512_ _0517_ VPWR VGND sg13g2_nand2_1
XFILLER_7_840 VPWR VGND sg13g2_decap_4
X_5880__389 VPWR VGND net389 sg13g2_tiehi
X_3461_ net542 net484 _0499_ VPWR VGND sg13g2_nor2_1
X_5200_ VGND VPWR _2033_ _2032_ _2031_ sg13g2_or2_1
X_3392_ VGND VPWR _0437_ _0438_ _0070_ _0439_ sg13g2_a21oi_1
X_5131_ _1970_ _1971_ _1972_ VPWR VGND sg13g2_nor2b_1
X_5062_ _1906_ mydesign.pe_weights\[32\] mydesign.pe_inputs\[22\] VPWR VGND sg13g2_nand2_1
X_4013_ _0973_ _0975_ _0987_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_917 VPWR VGND sg13g2_fill_1
XFILLER_41_909 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_17_clk clknet_3_3__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
X_5964_ net229 VGND VPWR net883 mydesign.accum\[74\] clknet_leaf_40_clk sg13g2_dfrbpq_2
X_4915_ net633 VPWR _1779_ VGND net1037 net442 sg13g2_o21ai_1
X_5895_ net363 VGND VPWR _0121_ mydesign.pe_weights\[53\] clknet_leaf_41_clk sg13g2_dfrbpq_2
X_4846_ net479 VPWR _1724_ VGND net582 net926 sg13g2_o21ai_1
X_4777_ _1658_ mydesign.accum\[49\] mydesign.pe_weights\[41\] net529 VPWR VGND sg13g2_and3_2
XFILLER_4_309 VPWR VGND sg13g2_decap_4
XFILLER_10_1019 VPWR VGND sg13g2_decap_8
X_3728_ VGND VPWR mydesign.accum\[116\] _0714_ _0737_ _0716_ sg13g2_a21oi_1
X_3659_ net480 VPWR _0672_ VGND net578 net851 sg13g2_o21ai_1
X_5329_ _2144_ VPWR _2146_ VGND _2142_ _2143_ sg13g2_o21ai_1
XFILLER_0_548 VPWR VGND sg13g2_decap_4
XFILLER_44_736 VPWR VGND sg13g2_decap_8
XFILLER_28_298 VPWR VGND sg13g2_decap_8
XFILLER_19_1011 VPWR VGND sg13g2_decap_8
XFILLER_40_931 VPWR VGND sg13g2_decap_8
XFILLER_25_994 VPWR VGND sg13g2_decap_8
X_5786__165 VPWR VGND net165 sg13g2_tiehi
XFILLER_21_8 VPWR VGND sg13g2_fill_1
XFILLER_19_298 VPWR VGND sg13g2_fill_2
XFILLER_35_725 VPWR VGND sg13g2_decap_4
XFILLER_22_408 VPWR VGND sg13g2_decap_8
X_5680_ _2464_ net645 _2461_ VPWR VGND sg13g2_nand2_1
XFILLER_31_964 VPWR VGND sg13g2_decap_8
X_4700_ VGND VPWR _1575_ _1583_ _1594_ _1582_ sg13g2_a21oi_1
XFILLER_33_1008 VPWR VGND sg13g2_decap_8
X_4631_ _1533_ VPWR _1534_ VGND net557 mydesign.inputs\[2\]\[11\] sg13g2_o21ai_1
XFILLER_30_496 VPWR VGND sg13g2_fill_1
X_4562_ _1451_ VPWR _1472_ VGND _1440_ _1452_ sg13g2_o21ai_1
X_4493_ net633 VPWR _1409_ VGND net530 net440 sg13g2_o21ai_1
X_3513_ net455 _0523_ mydesign.accum\[122\] _0541_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_6_clk clknet_3_1__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
X_3444_ _0405_ VPWR _0487_ VGND net509 _0484_ sg13g2_o21ai_1
XFILLER_40_0 VPWR VGND sg13g2_fill_2
X_3375_ VGND VPWR mydesign.accum\[9\] net514 _0424_ _0423_ sg13g2_a21oi_1
X_5114_ _1934_ VPWR _1956_ VGND _1923_ _1935_ sg13g2_o21ai_1
X_6094_ net324 VGND VPWR net417 mydesign.inputs\[3\]\[8\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_5045_ VGND VPWR _2530_ net442 _0270_ _1892_ sg13g2_a21oi_1
XFILLER_38_585 VPWR VGND sg13g2_fill_1
X_5947_ net263 VGND VPWR net984 mydesign.accum\[81\] clknet_leaf_25_clk sg13g2_dfrbpq_2
XFILLER_22_975 VPWR VGND sg13g2_decap_8
X_5878_ net393 VGND VPWR _0104_ mydesign.accum\[112\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_4829_ net533 mydesign.pe_inputs\[29\] mydesign.accum\[52\] _1707_ VPWR VGND sg13g2_nand3_1
XFILLER_1_857 VPWR VGND sg13g2_decap_4
XFILLER_49_839 VPWR VGND sg13g2_decap_8
XFILLER_1_1006 VPWR VGND sg13g2_decap_8
XFILLER_44_555 VPWR VGND sg13g2_decap_8
XFILLER_44_588 VPWR VGND sg13g2_fill_2
XFILLER_16_268 VPWR VGND sg13g2_fill_1
XFILLER_13_931 VPWR VGND sg13g2_decap_8
XFILLER_31_227 VPWR VGND sg13g2_fill_2
XFILLER_40_761 VPWR VGND sg13g2_fill_1
XFILLER_33_93 VPWR VGND sg13g2_fill_1
XFILLER_8_467 VPWR VGND sg13g2_decap_8
X_5879__391 VPWR VGND net391 sg13g2_tiehi
X_3160_ net499 net611 _2601_ VPWR VGND sg13g2_nor2_1
Xhold1 mydesign.cp2\[2\] VPWR VGND net407 sg13g2_dlygate4sd3_1
X_3091_ VPWR _2532_ net1033 VGND sg13g2_inv_1
XFILLER_23_706 VPWR VGND sg13g2_fill_1
X_5801_ net149 VGND VPWR _0027_ mydesign.inputs\[1\]\[14\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_23_739 VPWR VGND sg13g2_fill_2
X_3993_ _0968_ mydesign.pe_inputs\[53\] _0926_ VPWR VGND sg13g2_nand2_1
X_5732_ _2494_ VPWR _0355_ VGND net598 _2490_ sg13g2_o21ai_1
X_5663_ _2451_ _2444_ _2450_ VPWR VGND sg13g2_xnor2_1
X_5594_ net476 VPWR _2386_ VGND net586 net1040 sg13g2_o21ai_1
X_4614_ _0397_ _1518_ _1519_ _1520_ VPWR VGND sg13g2_nor3_1
X_4545_ _1455_ _1438_ _1456_ VPWR VGND sg13g2_nor2b_1
Xhold401 mydesign.accum\[18\] VPWR VGND net1020 sg13g2_dlygate4sd3_1
Xhold423 mydesign.accum\[20\] VPWR VGND net1042 sg13g2_dlygate4sd3_1
Xhold445 mydesign.load_counter\[3\] VPWR VGND net1064 sg13g2_dlygate4sd3_1
Xhold434 mydesign.accum\[96\] VPWR VGND net1053 sg13g2_dlygate4sd3_1
Xhold412 mydesign.pe_inputs\[26\] VPWR VGND net1031 sg13g2_dlygate4sd3_1
Xhold467 mydesign.pe_inputs\[62\] VPWR VGND net1086 sg13g2_dlygate4sd3_1
Xhold478 mydesign.pe_inputs\[20\] VPWR VGND net1097 sg13g2_dlygate4sd3_1
Xhold456 net12 VPWR VGND net1075 sg13g2_dlygate4sd3_1
X_4476_ net480 VPWR _1399_ VGND net581 net977 sg13g2_o21ai_1
Xhold489 mydesign.load_counter\[2\] VPWR VGND net1108 sg13g2_dlygate4sd3_1
X_3427_ net515 mydesign.accum\[110\] mydesign.accum\[78\] mydesign.accum\[46\] mydesign.accum\[14\]
+ net508 _0471_ VPWR VGND sg13g2_mux4_1
X_6146_ net164 VGND VPWR _0372_ mydesign.weights\[1\]\[20\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_3358_ net511 mydesign.accum\[120\] mydesign.accum\[88\] mydesign.accum\[56\] mydesign.accum\[24\]
+ net505 _0408_ VPWR VGND sg13g2_mux4_1
X_3289_ _2668_ net779 _2687_ _0042_ VPWR VGND sg13g2_mux2_1
X_6077_ net96 VGND VPWR _0303_ mydesign.accum\[19\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_5028_ _1865_ _1868_ _1879_ _1880_ VPWR VGND sg13g2_or3_1
XFILLER_26_533 VPWR VGND sg13g2_fill_2
XFILLER_9_209 VPWR VGND sg13g2_fill_2
XFILLER_10_923 VPWR VGND sg13g2_fill_1
XFILLER_6_927 VPWR VGND sg13g2_decap_4
XFILLER_10_956 VPWR VGND sg13g2_decap_8
XFILLER_5_448 VPWR VGND sg13g2_fill_1
X_5857__59 VPWR VGND net59 sg13g2_tiehi
XFILLER_0_142 VPWR VGND sg13g2_decap_8
XFILLER_0_153 VPWR VGND sg13g2_fill_1
XFILLER_49_636 VPWR VGND sg13g2_decap_8
X_5872__29 VPWR VGND net29 sg13g2_tiehi
XFILLER_17_511 VPWR VGND sg13g2_decap_4
XFILLER_29_360 VPWR VGND sg13g2_fill_1
XFILLER_45_842 VPWR VGND sg13g2_decap_8
XFILLER_17_544 VPWR VGND sg13g2_fill_2
XFILLER_44_396 VPWR VGND sg13g2_fill_2
XFILLER_32_525 VPWR VGND sg13g2_fill_2
XFILLER_13_794 VPWR VGND sg13g2_fill_2
XFILLER_8_253 VPWR VGND sg13g2_fill_2
X_4330_ _1252_ VPWR _1270_ VGND _1250_ _1253_ sg13g2_o21ai_1
XFILLER_5_993 VPWR VGND sg13g2_decap_8
X_4261_ _1205_ _1187_ _1204_ VPWR VGND sg13g2_nand2_1
XFILLER_4_481 VPWR VGND sg13g2_decap_4
X_6000_ net94 VGND VPWR _0226_ mydesign.accum\[62\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_3212_ _2606_ _2639_ _2640_ VPWR VGND sg13g2_nor2_2
X_4192_ _1149_ _1140_ _1148_ VPWR VGND sg13g2_nand2_1
X_3143_ VPWR _2584_ net407 VGND sg13g2_inv_1
XFILLER_36_842 VPWR VGND sg13g2_decap_8
X_3976_ _0926_ mydesign.pe_inputs\[52\] mydesign.accum\[98\] _0952_ VPWR VGND sg13g2_a21o_1
X_5925__307 VPWR VGND net307 sg13g2_tiehi
X_5715_ _2518_ _2484_ _2487_ VPWR VGND sg13g2_nor2_2
X_5646_ _2435_ _2430_ _2434_ VPWR VGND sg13g2_nand2_1
Xhold220 _0154_ VPWR VGND net839 sg13g2_dlygate4sd3_1
X_5577_ net749 mydesign.pe_inputs\[4\] net523 _2368_ _2370_ VPWR VGND sg13g2_and4_1
Xhold242 mydesign.accum\[69\] VPWR VGND net861 sg13g2_dlygate4sd3_1
Xhold253 mydesign.pe_weights\[49\] VPWR VGND net872 sg13g2_dlygate4sd3_1
X_4528_ _1430_ VPWR _1439_ VGND _1423_ _1431_ sg13g2_o21ai_1
Xhold231 _0253_ VPWR VGND net850 sg13g2_dlygate4sd3_1
Xhold275 mydesign.accum\[70\] VPWR VGND net894 sg13g2_dlygate4sd3_1
Xhold264 _0190_ VPWR VGND net883 sg13g2_dlygate4sd3_1
X_5901__351 VPWR VGND net351 sg13g2_tiehi
Xhold286 mydesign.accum\[77\] VPWR VGND net905 sg13g2_dlygate4sd3_1
X_4459_ mydesign.pe_inputs\[43\] net538 mydesign.accum\[78\] _1383_ VPWR VGND sg13g2_a21o_1
Xhold297 mydesign.accum\[105\] VPWR VGND net916 sg13g2_dlygate4sd3_1
XFILLER_18_308 VPWR VGND sg13g2_fill_2
X_6129_ net372 VGND VPWR net715 mydesign.weights\[0\]\[27\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_46_628 VPWR VGND sg13g2_decap_8
XFILLER_45_149 VPWR VGND sg13g2_fill_2
XFILLER_42_823 VPWR VGND sg13g2_fill_1
X_6016__26 VPWR VGND net26 sg13g2_tiehi
XFILLER_42_856 VPWR VGND sg13g2_decap_8
XFILLER_14_536 VPWR VGND sg13g2_decap_8
XFILLER_14_51 VPWR VGND sg13g2_fill_1
XFILLER_14_95 VPWR VGND sg13g2_fill_1
XFILLER_6_757 VPWR VGND sg13g2_fill_2
X_5976__205 VPWR VGND net205 sg13g2_tiehi
XFILLER_2_985 VPWR VGND sg13g2_decap_8
XFILLER_7_1023 VPWR VGND sg13g2_decap_4
XFILLER_37_606 VPWR VGND sg13g2_fill_2
XFILLER_49_499 VPWR VGND sg13g2_decap_8
XFILLER_44_160 VPWR VGND sg13g2_fill_2
XFILLER_32_311 VPWR VGND sg13g2_decap_8
X_3830_ _0822_ mydesign.pe_inputs\[57\] _0789_ VPWR VGND sg13g2_nand2_1
X_3761_ net471 VPWR _0768_ VGND net571 net973 sg13g2_o21ai_1
X_5500_ _2301_ _2298_ _2302_ VPWR VGND sg13g2_xor2_1
X_3692_ _0700_ _0701_ _0689_ _0703_ VPWR VGND sg13g2_nand3_1
X_5431_ _2242_ _2238_ _2241_ VPWR VGND sg13g2_xnor2_1
X_5362_ _2175_ _2154_ _2177_ VPWR VGND sg13g2_xor2_1
X_4313_ _1251_ _1253_ _1254_ VPWR VGND sg13g2_nor2_1
X_5293_ VGND VPWR _2094_ _2107_ _2121_ _2106_ sg13g2_a21oi_1
X_4244_ _1187_ _1188_ _1189_ VPWR VGND sg13g2_nor2b_1
X_4175_ VGND VPWR _1110_ _1112_ _1133_ _1132_ sg13g2_a21oi_1
X_3126_ _2567_ net995 VPWR VGND sg13g2_inv_2
XFILLER_35_28 VPWR VGND sg13g2_decap_4
XFILLER_24_834 VPWR VGND sg13g2_fill_2
XFILLER_24_845 VPWR VGND sg13g2_decap_4
XFILLER_23_344 VPWR VGND sg13g2_fill_2
XFILLER_23_355 VPWR VGND sg13g2_decap_8
X_6006__70 VPWR VGND net70 sg13g2_tiehi
X_3959_ _0936_ net1053 _0937_ VPWR VGND sg13g2_xor2_1
X_5629_ _2419_ _2409_ _2418_ VPWR VGND sg13g2_nand2_1
XFILLER_3_716 VPWR VGND sg13g2_fill_1
Xfanout541 net543 net541 VPWR VGND sg13g2_buf_8
Xfanout530 net938 net530 VPWR VGND sg13g2_buf_8
XFILLER_47_915 VPWR VGND sg13g2_decap_8
Xfanout574 net576 net574 VPWR VGND sg13g2_buf_8
Xfanout563 net595 net563 VPWR VGND sg13g2_buf_8
Xfanout552 net553 net552 VPWR VGND sg13g2_buf_2
XFILLER_46_403 VPWR VGND sg13g2_fill_2
Xfanout596 net1093 net596 VPWR VGND sg13g2_buf_8
Xfanout585 net589 net585 VPWR VGND sg13g2_buf_8
XFILLER_19_628 VPWR VGND sg13g2_fill_1
XFILLER_41_130 VPWR VGND sg13g2_fill_2
XFILLER_30_804 VPWR VGND sg13g2_fill_2
XFILLER_42_697 VPWR VGND sg13g2_decap_4
XFILLER_6_532 VPWR VGND sg13g2_fill_2
XFILLER_6_521 VPWR VGND sg13g2_fill_2
XFILLER_6_576 VPWR VGND sg13g2_decap_4
XFILLER_44_7 VPWR VGND sg13g2_fill_2
XFILLER_49_230 VPWR VGND sg13g2_decap_4
XFILLER_38_937 VPWR VGND sg13g2_decap_8
XFILLER_2_76 VPWR VGND sg13g2_fill_1
XFILLER_49_296 VPWR VGND sg13g2_decap_8
X_6050__258 VPWR VGND net258 sg13g2_tiehi
X_5980_ net197 VGND VPWR net874 mydesign.accum\[66\] clknet_leaf_45_clk sg13g2_dfrbpq_2
XFILLER_46_992 VPWR VGND sg13g2_decap_8
X_5841__87 VPWR VGND net87 sg13g2_tiehi
X_4931_ VGND VPWR mydesign.pe_weights\[37\] net528 _1788_ mydesign.accum\[41\] sg13g2_a21oi_1
XFILLER_17_182 VPWR VGND sg13g2_fill_1
XFILLER_18_694 VPWR VGND sg13g2_fill_1
X_4862_ _1739_ _1719_ _1722_ _1738_ VPWR VGND sg13g2_and3_1
XFILLER_21_804 VPWR VGND sg13g2_decap_8
X_3813_ net474 VPWR _0807_ VGND net688 _0806_ sg13g2_o21ai_1
XFILLER_21_815 VPWR VGND sg13g2_fill_2
XFILLER_33_675 VPWR VGND sg13g2_fill_1
XFILLER_33_686 VPWR VGND sg13g2_fill_1
XFILLER_33_697 VPWR VGND sg13g2_fill_1
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
XFILLER_32_185 VPWR VGND sg13g2_fill_1
X_4793_ _1669_ _1672_ _1673_ VPWR VGND sg13g2_nor2_1
X_3744_ _0752_ _0749_ _0750_ VPWR VGND sg13g2_xnor2_1
X_3675_ VGND VPWR net577 _0685_ _0106_ _0686_ sg13g2_a21oi_1
X_5414_ mydesign.pe_inputs\[15\] net527 mydesign.accum\[22\] _2226_ VPWR VGND sg13g2_nand3_1
XFILLER_0_708 VPWR VGND sg13g2_decap_8
XFILLER_0_719 VPWR VGND sg13g2_fill_1
X_5345_ _2158_ _2142_ _2161_ VPWR VGND sg13g2_xor2_1
X_5276_ _2105_ _2095_ _2103_ VPWR VGND sg13g2_xnor2_1
X_4227_ VGND VPWR _2568_ net438 _0167_ _1177_ sg13g2_a21oi_1
XFILLER_29_937 VPWR VGND sg13g2_decap_8
X_4158_ _1114_ _1116_ _1117_ VPWR VGND sg13g2_nor2_1
XFILLER_46_49 VPWR VGND sg13g2_decap_4
XFILLER_28_447 VPWR VGND sg13g2_fill_1
X_4089_ net626 VPWR _1057_ VGND net489 _1056_ sg13g2_o21ai_1
XFILLER_44_918 VPWR VGND sg13g2_decap_8
XFILLER_16_609 VPWR VGND sg13g2_fill_1
X_3109_ VPWR _2550_ net952 VGND sg13g2_inv_1
XFILLER_24_664 VPWR VGND sg13g2_decap_8
XFILLER_47_712 VPWR VGND sg13g2_decap_8
XFILLER_4_1004 VPWR VGND sg13g2_decap_8
XFILLER_19_403 VPWR VGND sg13g2_fill_1
XFILLER_19_436 VPWR VGND sg13g2_fill_2
XFILLER_47_789 VPWR VGND sg13g2_decap_8
XFILLER_46_266 VPWR VGND sg13g2_fill_1
XFILLER_28_970 VPWR VGND sg13g2_decap_8
XFILLER_35_929 VPWR VGND sg13g2_decap_8
XFILLER_43_984 VPWR VGND sg13g2_decap_8
XFILLER_15_675 VPWR VGND sg13g2_fill_2
XFILLER_6_384 VPWR VGND sg13g2_decap_4
X_6021__382 VPWR VGND net382 sg13g2_tiehi
X_3460_ net554 mydesign.inputs\[0\]\[24\] mydesign.inputs\[0\]\[20\] mydesign.inputs\[0\]\[16\]
+ mydesign.inputs\[0\]\[12\] net544 _0498_ VPWR VGND sg13g2_mux4_1
X_3391_ net622 VPWR _0439_ VGND net1087 net430 sg13g2_o21ai_1
X_5130_ _1948_ _1969_ _1945_ _1971_ VPWR VGND sg13g2_nand3_1
XFILLER_42_1010 VPWR VGND sg13g2_decap_8
X_5061_ VGND VPWR net584 _1904_ _0273_ _1905_ sg13g2_a21oi_1
XFILLER_28_2 VPWR VGND sg13g2_fill_1
X_4012_ VGND VPWR net564 _0985_ _0143_ _0986_ sg13g2_a21oi_1
X_5774__240 VPWR VGND net240 sg13g2_tiehi
XFILLER_37_222 VPWR VGND sg13g2_fill_2
XFILLER_37_211 VPWR VGND sg13g2_fill_2
XFILLER_37_233 VPWR VGND sg13g2_decap_8
X_5963_ net231 VGND VPWR net876 mydesign.accum\[73\] clknet_leaf_41_clk sg13g2_dfrbpq_2
X_4914_ VGND VPWR _2539_ net442 _0253_ _1778_ sg13g2_a21oi_1
X_5894_ net365 VGND VPWR _0120_ mydesign.pe_weights\[52\] clknet_leaf_40_clk sg13g2_dfrbpq_2
XFILLER_21_601 VPWR VGND sg13g2_decap_8
XFILLER_34_984 VPWR VGND sg13g2_decap_8
X_4845_ VGND VPWR _1721_ _1722_ _1723_ net502 sg13g2_a21oi_1
XFILLER_20_144 VPWR VGND sg13g2_fill_2
X_4776_ VGND VPWR net745 _1656_ _0236_ _1657_ sg13g2_a21oi_1
X_3727_ _0735_ _0732_ _0736_ VPWR VGND sg13g2_xor2_1
XFILLER_20_177 VPWR VGND sg13g2_fill_1
XFILLER_20_188 VPWR VGND sg13g2_fill_1
X_3658_ _0671_ _0669_ _0670_ VPWR VGND sg13g2_nand2_1
X_3589_ net468 VPWR _0614_ VGND net558 net1060 sg13g2_o21ai_1
X_5328_ _2142_ _2143_ _2144_ _2145_ VPWR VGND sg13g2_nor3_1
X_5259_ _2089_ _2077_ _2087_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_222 VPWR VGND sg13g2_decap_8
XFILLER_44_715 VPWR VGND sg13g2_decap_8
XFILLER_40_910 VPWR VGND sg13g2_decap_8
XFILLER_24_450 VPWR VGND sg13g2_decap_4
XFILLER_25_973 VPWR VGND sg13g2_decap_8
XFILLER_40_987 VPWR VGND sg13g2_decap_8
XFILLER_7_104 VPWR VGND sg13g2_fill_2
XFILLER_11_166 VPWR VGND sg13g2_fill_1
XFILLER_3_343 VPWR VGND sg13g2_fill_2
XFILLER_26_1016 VPWR VGND sg13g2_decap_8
XFILLER_26_1027 VPWR VGND sg13g2_fill_2
X_5834__101 VPWR VGND net101 sg13g2_tiehi
XFILLER_19_266 VPWR VGND sg13g2_fill_1
XFILLER_43_781 VPWR VGND sg13g2_decap_8
XFILLER_16_984 VPWR VGND sg13g2_decap_8
XFILLER_31_943 VPWR VGND sg13g2_decap_8
X_5984__189 VPWR VGND net189 sg13g2_tiehi
X_4630_ VGND VPWR net557 _2594_ _1533_ _0397_ sg13g2_a21oi_1
X_4561_ _1469_ _1470_ _1471_ VPWR VGND sg13g2_and2_1
X_3512_ _0540_ _0506_ _0517_ VPWR VGND sg13g2_nand2_1
X_4492_ VGND VPWR _2555_ net441 _0201_ _1408_ sg13g2_a21oi_1
X_3443_ VGND VPWR mydesign.accum\[23\] net516 _0486_ _0485_ sg13g2_a21oi_1
X_5113_ _1953_ _1954_ _1955_ VPWR VGND sg13g2_and2_1
X_3374_ net514 mydesign.accum\[41\] _0423_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_0 VPWR VGND sg13g2_decap_8
X_6093_ net332 VGND VPWR net1056 mydesign.accum\[15\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_5044_ net634 VPWR _1892_ VGND net1017 net443 sg13g2_o21ai_1
X_5946_ net265 VGND VPWR net740 mydesign.accum\[80\] clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_40_206 VPWR VGND sg13g2_decap_8
X_5877_ net395 VGND VPWR _0103_ mydesign.pe_weights\[59\] clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_22_954 VPWR VGND sg13g2_decap_8
X_4828_ _1706_ mydesign.pe_weights\[42\] mydesign.pe_inputs\[30\] VPWR VGND sg13g2_nand2_1
XFILLER_33_291 VPWR VGND sg13g2_fill_2
X_4759_ VGND VPWR _2547_ net450 _0228_ _1648_ sg13g2_a21oi_1
X_5869__35 VPWR VGND net35 sg13g2_tiehi
XFILLER_1_836 VPWR VGND sg13g2_decap_4
XFILLER_0_324 VPWR VGND sg13g2_decap_8
XFILLER_49_818 VPWR VGND sg13g2_decap_8
XFILLER_0_368 VPWR VGND sg13g2_fill_2
XFILLER_44_545 VPWR VGND sg13g2_fill_1
XFILLER_12_420 VPWR VGND sg13g2_decap_4
XFILLER_12_442 VPWR VGND sg13g2_fill_2
XFILLER_13_987 VPWR VGND sg13g2_decap_8
XFILLER_32_1020 VPWR VGND sg13g2_decap_8
X_3090_ VPWR _2531_ net828 VGND sg13g2_inv_1
XFILLER_0_880 VPWR VGND sg13g2_decap_8
Xhold2 _0067_ VPWR VGND net408 sg13g2_dlygate4sd3_1
XFILLER_48_895 VPWR VGND sg13g2_decap_8
XFILLER_35_512 VPWR VGND sg13g2_decap_4
X_5800_ net150 VGND VPWR _0026_ mydesign.inputs\[1\]\[13\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3992_ _0967_ mydesign.pe_inputs\[54\] _0919_ VPWR VGND sg13g2_nand2_1
XFILLER_16_792 VPWR VGND sg13g2_decap_4
X_5731_ net714 _2490_ net620 _2494_ VPWR VGND sg13g2_nand3_1
XFILLER_31_740 VPWR VGND sg13g2_fill_2
X_5662_ VPWR _2450_ _2449_ VGND sg13g2_inv_1
X_5593_ _2385_ _2370_ _2383_ VPWR VGND sg13g2_xnor2_1
X_4613_ mydesign.inputs\[2\]\[4\] net557 _1519_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_980 VPWR VGND sg13g2_decap_8
X_4544_ _1455_ _1439_ _1453_ VPWR VGND sg13g2_xnor2_1
Xhold402 _0302_ VPWR VGND net1021 sg13g2_dlygate4sd3_1
XFILLER_7_490 VPWR VGND sg13g2_fill_2
Xhold435 _0937_ VPWR VGND net1054 sg13g2_dlygate4sd3_1
Xhold424 mydesign.pe_weights\[20\] VPWR VGND net1043 sg13g2_dlygate4sd3_1
Xhold413 _0230_ VPWR VGND net1032 sg13g2_dlygate4sd3_1
Xhold457 mydesign.pe_inputs\[52\] VPWR VGND net1076 sg13g2_dlygate4sd3_1
Xhold446 mydesign.pe_inputs\[4\] VPWR VGND net1065 sg13g2_dlygate4sd3_1
Xhold468 net10 VPWR VGND net1087 sg13g2_dlygate4sd3_1
X_4475_ _1398_ _1394_ _1397_ VPWR VGND sg13g2_xnor2_1
X_3426_ VGND VPWR net456 _0469_ _0470_ _2698_ sg13g2_a21oi_1
Xhold479 mydesign.pe_inputs\[12\] VPWR VGND net1098 sg13g2_dlygate4sd3_1
X_3357_ net755 net834 _0407_ VPWR VGND sg13g2_nor2_1
X_6145_ net184 VGND VPWR _0371_ mydesign.weights\[0\]\[15\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5893__367 VPWR VGND net367 sg13g2_tiehi
X_6076_ net104 VGND VPWR net1021 mydesign.accum\[18\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_5027_ _1879_ _1871_ _1878_ VPWR VGND sg13g2_xnor2_1
X_3288_ _2667_ net795 _2687_ _0041_ VPWR VGND sg13g2_mux2_1
XFILLER_38_372 VPWR VGND sg13g2_fill_1
XFILLER_41_548 VPWR VGND sg13g2_fill_2
X_5929_ net299 VGND VPWR _0155_ mydesign.pe_weights\[47\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_16_1026 VPWR VGND sg13g2_fill_2
XFILLER_10_913 VPWR VGND sg13g2_fill_1
XFILLER_49_615 VPWR VGND sg13g2_decap_8
XFILLER_1_699 VPWR VGND sg13g2_fill_2
XFILLER_23_1008 VPWR VGND sg13g2_decap_8
X_6121__64 VPWR VGND net64 sg13g2_tiehi
XFILLER_45_821 VPWR VGND sg13g2_decap_8
XFILLER_28_61 VPWR VGND sg13g2_fill_1
XFILLER_45_898 VPWR VGND sg13g2_decap_8
XFILLER_44_342 VPWR VGND sg13g2_decap_8
XFILLER_44_82 VPWR VGND sg13g2_decap_8
XFILLER_9_711 VPWR VGND sg13g2_fill_1
X_6046__274 VPWR VGND net274 sg13g2_tiehi
XFILLER_5_972 VPWR VGND sg13g2_decap_8
X_4260_ _1204_ _1194_ _1203_ VPWR VGND sg13g2_xnor2_1
X_4191_ _1148_ _1145_ _1146_ VPWR VGND sg13g2_xnor2_1
X_3211_ _2639_ mydesign.load_counter\[3\] VPWR VGND net1108 sg13g2_nand2b_2
XFILLER_39_114 VPWR VGND sg13g2_decap_8
X_3142_ VPWR _2583_ net1073 VGND sg13g2_inv_1
XFILLER_48_692 VPWR VGND sg13g2_decap_8
XFILLER_39_1026 VPWR VGND sg13g2_fill_2
X_3975_ VPWR _0951_ _0950_ VGND sg13g2_inv_1
X_5714_ net774 _2486_ _2481_ _0345_ VPWR VGND sg13g2_mux2_1
X_5645_ _2433_ _2432_ _2434_ VPWR VGND sg13g2_xor2_1
X_6101__268 VPWR VGND net268 sg13g2_tiehi
Xhold210 _0269_ VPWR VGND net829 sg13g2_dlygate4sd3_1
X_5576_ mydesign.pe_inputs\[4\] net524 net749 _2369_ VPWR VGND sg13g2_nand3_1
Xhold221 mydesign.accum\[61\] VPWR VGND net840 sg13g2_dlygate4sd3_1
X_4527_ _1434_ VPWR _1438_ VGND _1420_ _1435_ sg13g2_o21ai_1
Xhold243 mydesign.pe_weights\[37\] VPWR VGND net862 sg13g2_dlygate4sd3_1
Xhold232 mydesign.accum\[113\] VPWR VGND net851 sg13g2_dlygate4sd3_1
Xhold276 mydesign.accum\[86\] VPWR VGND net895 sg13g2_dlygate4sd3_1
Xhold265 mydesign.accum\[62\] VPWR VGND net884 sg13g2_dlygate4sd3_1
Xhold287 mydesign.accum\[67\] VPWR VGND net906 sg13g2_dlygate4sd3_1
Xhold254 mydesign.accum\[66\] VPWR VGND net873 sg13g2_dlygate4sd3_1
X_4458_ net538 mydesign.pe_inputs\[43\] mydesign.accum\[78\] _1382_ VPWR VGND sg13g2_nand3_1
Xhold298 _0125_ VPWR VGND net917 sg13g2_dlygate4sd3_1
X_3409_ _0455_ _0454_ net457 _0452_ net456 VPWR VGND sg13g2_a22oi_1
X_4389_ _1314_ _1298_ _1317_ VPWR VGND sg13g2_xor2_1
X_6128_ net384 VGND VPWR _0354_ mydesign.weights\[0\]\[26\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_46_607 VPWR VGND sg13g2_decap_8
X_6059_ net222 VGND VPWR net955 mydesign.accum\[25\] clknet_leaf_6_clk sg13g2_dfrbpq_2
XFILLER_42_835 VPWR VGND sg13g2_decap_8
XFILLER_27_898 VPWR VGND sg13g2_decap_4
XFILLER_41_345 VPWR VGND sg13g2_decap_8
X_6145__184 VPWR VGND net184 sg13g2_tiehi
XFILLER_22_581 VPWR VGND sg13g2_fill_1
XFILLER_5_224 VPWR VGND sg13g2_fill_1
XFILLER_5_268 VPWR VGND sg13g2_fill_1
XFILLER_30_62 VPWR VGND sg13g2_fill_1
XFILLER_2_964 VPWR VGND sg13g2_decap_8
XFILLER_49_423 VPWR VGND sg13g2_fill_2
XFILLER_7_1002 VPWR VGND sg13g2_decap_8
XFILLER_49_434 VPWR VGND sg13g2_fill_1
XFILLER_39_71 VPWR VGND sg13g2_fill_2
X_5838__93 VPWR VGND net93 sg13g2_tiehi
XFILLER_17_342 VPWR VGND sg13g2_fill_2
XFILLER_18_865 VPWR VGND sg13g2_fill_1
XFILLER_45_695 VPWR VGND sg13g2_decap_8
X_3760_ _0767_ _0763_ _0766_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_518 VPWR VGND sg13g2_fill_2
X_5430_ _2241_ _2239_ _2240_ VPWR VGND sg13g2_xnor2_1
X_3691_ _0702_ _0689_ _0700_ _0701_ VPWR VGND sg13g2_and3_1
X_5361_ _2154_ _2175_ _2176_ VPWR VGND sg13g2_nor2b_1
X_4312_ VGND VPWR mydesign.pe_weights\[59\] mydesign.pe_inputs\[46\] _1253_ mydesign.accum\[85\]
+ sg13g2_a21oi_1
X_5292_ _2120_ _2104_ _2118_ VPWR VGND sg13g2_xnor2_1
X_4243_ _1186_ VPWR _1188_ VGND _1184_ _1185_ sg13g2_o21ai_1
X_6135__320 VPWR VGND net320 sg13g2_tiehi
X_4174_ _1130_ _1120_ _1132_ VPWR VGND sg13g2_xor2_1
X_3125_ VPWR _2566_ net989 VGND sg13g2_inv_1
XFILLER_35_150 VPWR VGND sg13g2_decap_8
XFILLER_24_868 VPWR VGND sg13g2_fill_2
XFILLER_23_367 VPWR VGND sg13g2_decap_8
XFILLER_23_378 VPWR VGND sg13g2_fill_1
X_3958_ _0936_ net564 _0935_ VPWR VGND sg13g2_nand2_1
X_3889_ mydesign.pe_inputs\[58\] _0804_ _0878_ VPWR VGND sg13g2_and2_1
X_5628_ _2418_ _2410_ _2416_ VPWR VGND sg13g2_xnor2_1
X_5559_ _2357_ net416 _2356_ VPWR VGND sg13g2_nand2_1
Xfanout531 net1101 net531 VPWR VGND sg13g2_buf_2
Xfanout520 mydesign.pe_inputs\[11\] net520 VPWR VGND sg13g2_buf_8
Xfanout542 net543 net542 VPWR VGND sg13g2_buf_8
Xfanout553 mydesign.cp\[0\] net553 VPWR VGND sg13g2_buf_8
Xfanout575 net576 net575 VPWR VGND sg13g2_buf_8
Xfanout564 net565 net564 VPWR VGND sg13g2_buf_8
Xfanout586 net587 net586 VPWR VGND sg13g2_buf_8
XFILLER_18_106 VPWR VGND sg13g2_fill_1
Xfanout597 _2631_ net597 VPWR VGND sg13g2_buf_8
XFILLER_27_651 VPWR VGND sg13g2_decap_8
XFILLER_15_846 VPWR VGND sg13g2_fill_2
XFILLER_30_827 VPWR VGND sg13g2_fill_2
XFILLER_41_197 VPWR VGND sg13g2_fill_1
XFILLER_23_890 VPWR VGND sg13g2_decap_8
XFILLER_41_61 VPWR VGND sg13g2_fill_1
XFILLER_29_1014 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_fill_2
XFILLER_1_282 VPWR VGND sg13g2_fill_1
XFILLER_38_916 VPWR VGND sg13g2_decap_8
XFILLER_37_415 VPWR VGND sg13g2_fill_2
XFILLER_37_426 VPWR VGND sg13g2_fill_1
XFILLER_46_971 VPWR VGND sg13g2_decap_8
X_4930_ _1787_ mydesign.accum\[41\] mydesign.pe_weights\[37\] net528 VPWR VGND sg13g2_and3_2
XFILLER_33_610 VPWR VGND sg13g2_decap_4
X_4861_ _1738_ _1715_ _1736_ VPWR VGND sg13g2_xnor2_1
XFILLER_17_194 VPWR VGND sg13g2_fill_1
XFILLER_36_1007 VPWR VGND sg13g2_decap_8
X_3812_ _0806_ net572 mydesign.pe_inputs\[56\] _0783_ VPWR VGND sg13g2_and3_1
XFILLER_20_304 VPWR VGND sg13g2_decap_8
X_4792_ _1672_ _1670_ _1671_ VPWR VGND sg13g2_nand2_1
X_3743_ VPWR _0751_ _0750_ VGND sg13g2_inv_1
XFILLER_9_360 VPWR VGND sg13g2_fill_2
X_3674_ net470 VPWR _0686_ VGND net577 net877 sg13g2_o21ai_1
X_5413_ _2225_ _2224_ _0305_ VPWR VGND sg13g2_nor2b_1
X_5344_ _2142_ _2158_ _2160_ VPWR VGND sg13g2_nor2_1
X_5275_ _2104_ _2095_ _2103_ VPWR VGND sg13g2_nand2_1
X_4226_ net630 VPWR _1177_ VGND mydesign.pe_inputs\[43\] net438 sg13g2_o21ai_1
X_4157_ VGND VPWR _1112_ _1113_ _1116_ _1097_ sg13g2_a21oi_1
XFILLER_29_916 VPWR VGND sg13g2_decap_8
XFILLER_28_437 VPWR VGND sg13g2_fill_1
X_3108_ VPWR _2549_ net535 VGND sg13g2_inv_1
X_4088_ _0639_ net791 _1055_ _1056_ VPWR VGND sg13g2_a21o_2
XFILLER_43_429 VPWR VGND sg13g2_decap_4
XFILLER_12_805 VPWR VGND sg13g2_fill_1
XFILLER_11_53 VPWR VGND sg13g2_decap_4
XFILLER_47_768 VPWR VGND sg13g2_decap_8
XFILLER_35_908 VPWR VGND sg13g2_decap_8
XFILLER_43_963 VPWR VGND sg13g2_decap_8
XFILLER_15_654 VPWR VGND sg13g2_fill_2
XFILLER_15_687 VPWR VGND sg13g2_decap_8
XFILLER_30_679 VPWR VGND sg13g2_fill_1
XFILLER_10_370 VPWR VGND sg13g2_fill_1
X_3390_ VPWR VGND net456 _0436_ _0430_ _0412_ _0438_ _0429_ sg13g2_a221oi_1
X_5060_ net475 VPWR _1905_ VGND net584 net919 sg13g2_o21ai_1
XFILLER_38_713 VPWR VGND sg13g2_fill_2
X_4011_ net466 VPWR _0986_ VGND net564 net967 sg13g2_o21ai_1
XFILLER_38_735 VPWR VGND sg13g2_fill_2
X_5962_ net233 VGND VPWR net685 mydesign.accum\[72\] clknet_leaf_40_clk sg13g2_dfrbpq_2
XFILLER_37_267 VPWR VGND sg13g2_fill_1
X_4913_ net634 VPWR _1778_ VGND mydesign.pe_inputs\[21\] net442 sg13g2_o21ai_1
XFILLER_34_963 VPWR VGND sg13g2_decap_8
X_5893_ net367 VGND VPWR net1047 mydesign.pe_inputs\[55\] clknet_leaf_43_clk sg13g2_dfrbpq_2
XFILLER_21_613 VPWR VGND sg13g2_fill_2
XFILLER_20_123 VPWR VGND sg13g2_decap_8
XFILLER_33_495 VPWR VGND sg13g2_decap_8
X_4844_ _1720_ VPWR _1722_ VGND _1699_ _1701_ sg13g2_o21ai_1
X_4775_ net480 VPWR _1657_ VGND net745 _1656_ sg13g2_o21ai_1
X_3726_ _0735_ _0733_ _0734_ VPWR VGND sg13g2_nand2_1
X_3657_ _0660_ mydesign.accum\[112\] _0668_ _0670_ VPWR VGND sg13g2_a21o_1
X_3588_ _0611_ _0598_ _0613_ VPWR VGND sg13g2_xor2_1
XFILLER_0_528 VPWR VGND sg13g2_decap_8
X_5327_ _2144_ mydesign.pe_inputs\[13\] mydesign.pe_weights\[24\] VPWR VGND sg13g2_nand2_1
X_5258_ _2088_ _2077_ _2087_ VPWR VGND sg13g2_nand2_1
X_4209_ VGND VPWR _1139_ _1152_ _1165_ _1151_ sg13g2_a21oi_1
X_5189_ _2023_ net563 _2022_ VPWR VGND sg13g2_nand2_1
XFILLER_43_215 VPWR VGND sg13g2_fill_2
XFILLER_37_790 VPWR VGND sg13g2_fill_2
XFILLER_25_952 VPWR VGND sg13g2_decap_8
XFILLER_40_966 VPWR VGND sg13g2_decap_8
XFILLER_4_867 VPWR VGND sg13g2_fill_1
XFILLER_3_377 VPWR VGND sg13g2_fill_1
XFILLER_47_565 VPWR VGND sg13g2_fill_2
XFILLER_43_760 VPWR VGND sg13g2_decap_8
XFILLER_16_963 VPWR VGND sg13g2_decap_8
XFILLER_31_922 VPWR VGND sg13g2_decap_8
X_4560_ _1447_ _1449_ _1468_ _1470_ VPWR VGND sg13g2_or3_1
XFILLER_31_999 VPWR VGND sg13g2_decap_8
X_4491_ net633 VPWR _1408_ VGND net828 net440 sg13g2_o21ai_1
X_3511_ VGND VPWR net558 _0538_ _0089_ _0539_ sg13g2_a21oi_1
X_3442_ net516 mydesign.accum\[55\] _0485_ VPWR VGND sg13g2_nor2b_1
XFILLER_40_2 VPWR VGND sg13g2_fill_1
X_3373_ mydesign.accum\[105\] mydesign.accum\[73\] net514 _0422_ VPWR VGND sg13g2_mux2_1
X_5112_ _1930_ _1932_ _1952_ _1954_ VPWR VGND sg13g2_or3_1
X_6092_ net344 VGND VPWR _0318_ mydesign.accum\[14\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_5043_ VGND VPWR _2531_ net443 _0269_ _1891_ sg13g2_a21oi_1
XFILLER_26_705 VPWR VGND sg13g2_decap_8
XFILLER_25_248 VPWR VGND sg13g2_decap_8
X_5945_ net267 VGND VPWR _0171_ mydesign.pe_weights\[43\] clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_34_771 VPWR VGND sg13g2_decap_8
X_5876_ net397 VGND VPWR _0102_ mydesign.pe_weights\[58\] clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_22_933 VPWR VGND sg13g2_decap_8
XFILLER_33_270 VPWR VGND sg13g2_decap_4
X_4827_ _1688_ VPWR _1705_ VGND _1687_ _1690_ sg13g2_o21ai_1
X_6104__244 VPWR VGND net244 sg13g2_tiehi
X_4758_ net637 VPWR _1648_ VGND net1022 net450 sg13g2_o21ai_1
X_4689_ _1584_ _1574_ _1583_ VPWR VGND sg13g2_xnor2_1
X_3709_ _0719_ _0712_ _0717_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_303 VPWR VGND sg13g2_decap_8
XFILLER_1_815 VPWR VGND sg13g2_fill_2
X_6118__92 VPWR VGND net92 sg13g2_tiehi
XFILLER_0_336 VPWR VGND sg13g2_fill_2
XFILLER_48_329 VPWR VGND sg13g2_fill_1
X_6111__204 VPWR VGND net204 sg13g2_tiehi
XFILLER_17_705 VPWR VGND sg13g2_decap_8
XFILLER_32_708 VPWR VGND sg13g2_decap_8
XFILLER_9_926 VPWR VGND sg13g2_decap_8
XFILLER_13_966 VPWR VGND sg13g2_decap_8
XFILLER_4_653 VPWR VGND sg13g2_fill_2
XFILLER_4_631 VPWR VGND sg13g2_fill_1
XFILLER_4_675 VPWR VGND sg13g2_decap_4
X_6124__40 VPWR VGND net40 sg13g2_tiehi
Xhold3 mydesign.accum\[7\] VPWR VGND net409 sg13g2_dlygate4sd3_1
XFILLER_48_874 VPWR VGND sg13g2_decap_8
XFILLER_35_535 VPWR VGND sg13g2_fill_1
X_3991_ VPWR _0966_ _0965_ VGND sg13g2_inv_1
X_5730_ _2493_ VPWR _0354_ VGND net600 _2490_ sg13g2_o21ai_1
X_5661_ VGND VPWR _2449_ _2448_ _2447_ sg13g2_or2_1
X_5592_ _2384_ _2370_ _2383_ VPWR VGND sg13g2_nand2_1
X_4612_ net557 mydesign.inputs\[2\]\[8\] _1518_ VPWR VGND sg13g2_nor2_1
X_4543_ _1439_ _1453_ _1454_ VPWR VGND sg13g2_and2_1
Xhold425 mydesign.load_counter\[1\] VPWR VGND net1044 sg13g2_dlygate4sd3_1
Xhold414 mydesign.pe_weights\[32\] VPWR VGND net1033 sg13g2_dlygate4sd3_1
Xhold436 mydesign.accum\[15\] VPWR VGND net1055 sg13g2_dlygate4sd3_1
Xhold403 mydesign.pe_inputs\[24\] VPWR VGND net1022 sg13g2_dlygate4sd3_1
Xhold469 mydesign.cp\[1\] VPWR VGND net1088 sg13g2_dlygate4sd3_1
Xhold447 _0308_ VPWR VGND net1066 sg13g2_dlygate4sd3_1
X_4474_ _1397_ _1395_ _1396_ VPWR VGND sg13g2_xnor2_1
Xhold458 mydesign.pe_weights\[31\] VPWR VGND net1077 sg13g2_dlygate4sd3_1
X_3425_ net511 mydesign.accum\[126\] mydesign.accum\[94\] mydesign.accum\[62\] mydesign.accum\[30\]
+ net505 _0469_ VPWR VGND sg13g2_mux4_1
X_6144_ net200 VGND VPWR _0370_ mydesign.weights\[0\]\[14\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3356_ net515 mydesign.accum\[112\] mydesign.accum\[80\] mydesign.accum\[48\] mydesign.accum\[16\]
+ net509 _0406_ VPWR VGND sg13g2_mux4_1
X_3287_ _2687_ _2655_ _2686_ VPWR VGND sg13g2_nand2_2
X_6075_ net112 VGND VPWR net1030 mydesign.accum\[17\] clknet_leaf_27_clk sg13g2_dfrbpq_2
XFILLER_39_841 VPWR VGND sg13g2_fill_2
X_5026_ _1878_ _1877_ _1876_ VPWR VGND sg13g2_nand2b_1
XFILLER_26_513 VPWR VGND sg13g2_decap_8
XFILLER_26_524 VPWR VGND sg13g2_fill_1
XFILLER_26_579 VPWR VGND sg13g2_decap_8
X_5928_ net301 VGND VPWR net839 mydesign.pe_weights\[46\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_16_1005 VPWR VGND sg13g2_decap_8
X_5859_ net55 VGND VPWR _0085_ mydesign.pe_weights\[61\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_21_251 VPWR VGND sg13g2_fill_1
XFILLER_22_785 VPWR VGND sg13g2_decap_8
XFILLER_5_406 VPWR VGND sg13g2_fill_1
XFILLER_1_667 VPWR VGND sg13g2_fill_2
XFILLER_45_800 VPWR VGND sg13g2_decap_8
XFILLER_44_310 VPWR VGND sg13g2_fill_1
XFILLER_17_546 VPWR VGND sg13g2_fill_1
XFILLER_29_384 VPWR VGND sg13g2_fill_2
XFILLER_45_877 VPWR VGND sg13g2_decap_8
XFILLER_32_527 VPWR VGND sg13g2_fill_1
XFILLER_8_200 VPWR VGND sg13g2_fill_2
XFILLER_40_593 VPWR VGND sg13g2_fill_1
XFILLER_8_255 VPWR VGND sg13g2_fill_1
XFILLER_12_284 VPWR VGND sg13g2_fill_2
X_4190_ _1147_ _1145_ _1146_ VPWR VGND sg13g2_nand2b_1
X_3210_ _2588_ net596 _2638_ VPWR VGND sg13g2_nor2_1
X_5856__61 VPWR VGND net61 sg13g2_tiehi
X_6053__246 VPWR VGND net246 sg13g2_tiehi
X_3141_ VPWR _2582_ net1015 VGND sg13g2_inv_1
XFILLER_39_148 VPWR VGND sg13g2_fill_2
X_5871__31 VPWR VGND net31 sg13g2_tiehi
XFILLER_48_671 VPWR VGND sg13g2_decap_8
XFILLER_36_811 VPWR VGND sg13g2_fill_2
XFILLER_36_822 VPWR VGND sg13g2_fill_2
XFILLER_39_1005 VPWR VGND sg13g2_decap_8
X_3974_ mydesign.pe_inputs\[52\] _0926_ mydesign.accum\[98\] _0950_ VPWR VGND sg13g2_nand3_1
X_5713_ _2519_ _2484_ _2486_ VPWR VGND sg13g2_nor2_2
X_5644_ _2433_ net519 mydesign.pe_weights\[18\] VPWR VGND sg13g2_nand2_1
X_5575_ _2368_ _2363_ _2367_ VPWR VGND sg13g2_xnor2_1
Xhold211 mydesign.pe_weights\[38\] VPWR VGND net830 sg13g2_dlygate4sd3_1
Xhold200 _0221_ VPWR VGND net819 sg13g2_dlygate4sd3_1
Xhold222 mydesign.accum\[68\] VPWR VGND net841 sg13g2_dlygate4sd3_1
X_4526_ VGND VPWR net566 _1436_ _0206_ _1437_ sg13g2_a21oi_1
Xhold244 _0257_ VPWR VGND net863 sg13g2_dlygate4sd3_1
Xhold233 _0105_ VPWR VGND net852 sg13g2_dlygate4sd3_1
Xhold277 mydesign.accum\[89\] VPWR VGND net896 sg13g2_dlygate4sd3_1
XFILLER_49_28 VPWR VGND sg13g2_decap_8
Xhold255 _0206_ VPWR VGND net874 sg13g2_dlygate4sd3_1
Xhold266 mydesign.weights\[2\]\[15\] VPWR VGND net885 sg13g2_dlygate4sd3_1
X_4457_ net463 _1381_ _0193_ VPWR VGND sg13g2_nor2_1
Xhold299 mydesign.accum\[53\] VPWR VGND net918 sg13g2_dlygate4sd3_1
Xhold288 mydesign.accum\[65\] VPWR VGND net907 sg13g2_dlygate4sd3_1
X_3408_ net512 mydesign.accum\[100\] mydesign.accum\[68\] mydesign.accum\[36\] mydesign.accum\[4\]
+ net507 _0454_ VPWR VGND sg13g2_mux4_1
X_4388_ _1298_ _1314_ _1316_ VPWR VGND sg13g2_nor2_1
X_6127_ net392 VGND VPWR _0353_ mydesign.weights\[0\]\[25\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3339_ _0393_ net546 VPWR VGND net543 sg13g2_nand2b_2
X_6058_ net226 VGND VPWR _0284_ mydesign.accum\[24\] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_5009_ _1861_ VPWR _1862_ VGND _1840_ _1842_ sg13g2_o21ai_1
XFILLER_26_310 VPWR VGND sg13g2_fill_1
XFILLER_26_321 VPWR VGND sg13g2_fill_2
XFILLER_14_505 VPWR VGND sg13g2_fill_1
XFILLER_26_343 VPWR VGND sg13g2_decap_8
XFILLER_26_354 VPWR VGND sg13g2_fill_1
XFILLER_41_335 VPWR VGND sg13g2_fill_2
XFILLER_14_549 VPWR VGND sg13g2_fill_1
XFILLER_5_203 VPWR VGND sg13g2_fill_2
XFILLER_2_921 VPWR VGND sg13g2_fill_2
XFILLER_17_321 VPWR VGND sg13g2_decap_8
XFILLER_18_855 VPWR VGND sg13g2_fill_2
XFILLER_45_674 VPWR VGND sg13g2_decap_8
XFILLER_44_162 VPWR VGND sg13g2_fill_1
XFILLER_9_531 VPWR VGND sg13g2_fill_1
X_3690_ _0699_ _0698_ _0678_ _0701_ VPWR VGND sg13g2_a21o_1
X_5360_ _2174_ _2171_ _2175_ VPWR VGND sg13g2_xor2_1
X_4311_ mydesign.pe_weights\[59\] mydesign.pe_inputs\[46\] mydesign.accum\[85\] _1252_
+ VPWR VGND sg13g2_nand3_1
X_6094__324 VPWR VGND net324 sg13g2_tiehi
X_5291_ _2104_ _2118_ _2119_ VPWR VGND sg13g2_nor2b_1
X_4242_ _1184_ _1185_ _1186_ _1187_ VPWR VGND sg13g2_nor3_1
X_4173_ _1131_ _1130_ _1120_ VPWR VGND sg13g2_nand2b_1
X_3124_ VPWR _2565_ net988 VGND sg13g2_inv_1
XFILLER_27_129 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_47_clk clknet_3_1__leaf_clk clknet_leaf_47_clk VPWR VGND sg13g2_buf_8
XFILLER_23_313 VPWR VGND sg13g2_decap_4
XFILLER_36_674 VPWR VGND sg13g2_fill_2
XFILLER_23_346 VPWR VGND sg13g2_fill_1
XFILLER_35_184 VPWR VGND sg13g2_fill_1
X_3957_ _0914_ mydesign.pe_inputs\[52\] _0935_ VPWR VGND sg13g2_nor2b_1
XFILLER_13_1008 VPWR VGND sg13g2_decap_8
X_3888_ _0877_ mydesign.pe_inputs\[59\] _0796_ VPWR VGND sg13g2_nand2_1
X_5627_ _2417_ _2416_ _2410_ VPWR VGND sg13g2_nand2b_1
X_5558_ VGND VPWR net608 _2356_ _2354_ net606 sg13g2_a21oi_2
X_4509_ net473 VPWR _1422_ VGND net574 net907 sg13g2_o21ai_1
X_5489_ _2292_ _2276_ _2290_ VPWR VGND sg13g2_xnor2_1
Xfanout532 net1095 net532 VPWR VGND sg13g2_buf_8
Xfanout510 net1103 net510 VPWR VGND sg13g2_buf_8
Xfanout521 mydesign.pe_inputs\[8\] net521 VPWR VGND sg13g2_buf_8
Xfanout565 net566 net565 VPWR VGND sg13g2_buf_8
Xfanout543 net1083 net543 VPWR VGND sg13g2_buf_8
Xfanout554 net556 net554 VPWR VGND sg13g2_buf_8
Xfanout587 net588 net587 VPWR VGND sg13g2_buf_8
Xfanout576 net594 net576 VPWR VGND sg13g2_buf_8
Xfanout598 _2631_ net598 VPWR VGND sg13g2_buf_8
XFILLER_46_427 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_38_clk clknet_3_5__leaf_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_26_195 VPWR VGND sg13g2_fill_2
XFILLER_41_165 VPWR VGND sg13g2_fill_1
XFILLER_30_806 VPWR VGND sg13g2_fill_1
X_6012__42 VPWR VGND net42 sg13g2_tiehi
XFILLER_6_523 VPWR VGND sg13g2_fill_1
XFILLER_46_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_29_clk clknet_3_7__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_17_140 VPWR VGND sg13g2_fill_1
X_4860_ _1715_ _1736_ _1737_ VPWR VGND sg13g2_nor2_1
X_3811_ VGND VPWR _2556_ net492 _0123_ _0805_ sg13g2_a21oi_1
XFILLER_20_338 VPWR VGND sg13g2_fill_2
X_4791_ net529 mydesign.pe_weights\[42\] mydesign.accum\[50\] _1671_ VPWR VGND sg13g2_a21o_1
X_3742_ _0733_ VPWR _0750_ VGND _0732_ _0735_ sg13g2_o21ai_1
X_3673_ _0685_ _0669_ _0684_ VPWR VGND sg13g2_xnor2_1
X_5412_ net482 VPWR _2225_ VGND net590 net1035 sg13g2_o21ai_1
X_5343_ _2159_ _2142_ _2158_ VPWR VGND sg13g2_nand2_1
X_5274_ _2103_ _2100_ _2101_ VPWR VGND sg13g2_xnor2_1
X_4225_ VGND VPWR _2569_ net439 _0166_ _1176_ sg13g2_a21oi_1
X_4156_ _1112_ _1113_ _1097_ _1115_ VPWR VGND sg13g2_nand3_1
X_3107_ VPWR _2548_ mydesign.accum\[61\] VGND sg13g2_inv_1
X_4087_ VGND VPWR _1053_ _1054_ _1055_ net542 sg13g2_a21oi_1
XFILLER_37_994 VPWR VGND sg13g2_decap_8
XFILLER_36_471 VPWR VGND sg13g2_fill_1
X_4989_ _1841_ _1833_ _1843_ VPWR VGND sg13g2_xor2_1
XFILLER_3_526 VPWR VGND sg13g2_fill_1
XFILLER_11_98 VPWR VGND sg13g2_decap_8
XFILLER_47_747 VPWR VGND sg13g2_decap_8
XFILLER_43_942 VPWR VGND sg13g2_decap_8
XFILLER_42_430 VPWR VGND sg13g2_fill_1
XFILLER_14_110 VPWR VGND sg13g2_fill_2
XFILLER_14_154 VPWR VGND sg13g2_fill_2
XFILLER_15_677 VPWR VGND sg13g2_fill_1
XFILLER_35_5 VPWR VGND sg13g2_decap_4
X_4010_ _0985_ _0963_ _0984_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_460 VPWR VGND sg13g2_fill_2
XFILLER_19_983 VPWR VGND sg13g2_decap_8
X_5961_ net235 VGND VPWR _0187_ mydesign.pe_weights\[39\] clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_37_279 VPWR VGND sg13g2_fill_2
XFILLER_45_290 VPWR VGND sg13g2_decap_8
X_4912_ VGND VPWR _2540_ net442 _0252_ _1777_ sg13g2_a21oi_1
XFILLER_18_493 VPWR VGND sg13g2_decap_8
XFILLER_34_942 VPWR VGND sg13g2_decap_8
X_5892_ net369 VGND VPWR _0118_ mydesign.pe_inputs\[54\] clknet_leaf_43_clk sg13g2_dfrbpq_2
XFILLER_33_485 VPWR VGND sg13g2_decap_4
X_4843_ _1699_ _1701_ _1720_ _1721_ VPWR VGND sg13g2_or3_1
X_4774_ net502 _2544_ _2547_ _1656_ VPWR VGND sg13g2_nor3_1
X_3725_ _0658_ mydesign.pe_inputs\[62\] mydesign.accum\[117\] _0734_ VPWR VGND sg13g2_a21o_1
Xclkbuf_leaf_9_clk clknet_3_0__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_3656_ _0660_ _0668_ mydesign.accum\[112\] _0669_ VPWR VGND sg13g2_nand3_1
X_3587_ VGND VPWR _0592_ _0595_ _0612_ _0611_ sg13g2_a21oi_1
X_5326_ VGND VPWR net522 mydesign.pe_weights\[25\] _2143_ mydesign.accum\[17\] sg13g2_a21oi_1
X_5257_ _2086_ _2078_ _2087_ VPWR VGND sg13g2_xor2_1
X_5779__175 VPWR VGND net175 sg13g2_tiehi
X_4208_ _1164_ _1160_ _1163_ VPWR VGND sg13g2_xnor2_1
X_5188_ net891 _2004_ _2022_ VPWR VGND sg13g2_and2_1
X_4139_ _1098_ mydesign.pe_weights\[60\] _1061_ VPWR VGND sg13g2_nand2_1
XFILLER_28_246 VPWR VGND sg13g2_fill_1
XFILLER_19_1025 VPWR VGND sg13g2_decap_4
XFILLER_36_290 VPWR VGND sg13g2_fill_2
XFILLER_40_945 VPWR VGND sg13g2_decap_8
XFILLER_8_607 VPWR VGND sg13g2_fill_1
XFILLER_3_345 VPWR VGND sg13g2_fill_1
X_6090__360 VPWR VGND net360 sg13g2_tiehi
XFILLER_16_942 VPWR VGND sg13g2_decap_8
XFILLER_34_249 VPWR VGND sg13g2_decap_4
X_6049__262 VPWR VGND net262 sg13g2_tiehi
XFILLER_31_901 VPWR VGND sg13g2_decap_8
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_15_474 VPWR VGND sg13g2_decap_8
XFILLER_31_978 VPWR VGND sg13g2_decap_8
X_3510_ net467 VPWR _0539_ VGND net558 net937 sg13g2_o21ai_1
X_4490_ VGND VPWR _2532_ net493 _0200_ _1407_ sg13g2_a21oi_1
X_3441_ mydesign.accum\[119\] mydesign.accum\[87\] net516 _0484_ VPWR VGND sg13g2_mux2_1
X_3372_ net511 mydesign.accum\[121\] mydesign.accum\[89\] mydesign.accum\[57\] mydesign.accum\[25\]
+ net505 _0421_ VPWR VGND sg13g2_mux4_1
X_5111_ _1952_ VPWR _1953_ VGND _1930_ _1932_ sg13g2_o21ai_1
X_6091_ net352 VGND VPWR _0317_ mydesign.accum\[13\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_5042_ net634 VPWR _1891_ VGND mydesign.pe_weights\[17\] net443 sg13g2_o21ai_1
XFILLER_19_0 VPWR VGND sg13g2_fill_2
X_5932__293 VPWR VGND net293 sg13g2_tiehi
X_5944_ net269 VGND VPWR _0170_ mydesign.pe_weights\[42\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_5875_ net23 VGND VPWR _0101_ mydesign.pe_weights\[57\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4826_ _1704_ mydesign.pe_weights\[41\] mydesign.pe_inputs\[31\] VPWR VGND sg13g2_nand2_1
XFILLER_33_282 VPWR VGND sg13g2_fill_2
XFILLER_22_989 VPWR VGND sg13g2_decap_8
X_4757_ VGND VPWR net568 _1646_ _0227_ _1647_ sg13g2_a21oi_1
XFILLER_49_1007 VPWR VGND sg13g2_decap_8
X_4688_ _1583_ _1557_ _1581_ VPWR VGND sg13g2_xnor2_1
X_3708_ _0718_ _0712_ _0717_ VPWR VGND sg13g2_nand2_1
X_3639_ VGND VPWR _2565_ net492 _0102_ _0654_ sg13g2_a21oi_1
X_5309_ _2133_ VPWR _0293_ VGND net601 _2130_ sg13g2_o21ai_1
XFILLER_29_544 VPWR VGND sg13g2_decap_8
XFILLER_17_739 VPWR VGND sg13g2_fill_1
XFILLER_29_599 VPWR VGND sg13g2_fill_2
XFILLER_44_569 VPWR VGND sg13g2_decap_4
XFILLER_13_901 VPWR VGND sg13g2_fill_2
XFILLER_17_75 VPWR VGND sg13g2_decap_8
XFILLER_17_86 VPWR VGND sg13g2_fill_1
XFILLER_13_945 VPWR VGND sg13g2_decap_8
XFILLER_12_444 VPWR VGND sg13g2_fill_1
XFILLER_33_52 VPWR VGND sg13g2_decap_8
XFILLER_40_797 VPWR VGND sg13g2_fill_2
XFILLER_8_426 VPWR VGND sg13g2_fill_1
X_5983__191 VPWR VGND net191 sg13g2_tiehi
XFILLER_12_466 VPWR VGND sg13g2_decap_8
XFILLER_4_643 VPWR VGND sg13g2_fill_2
XFILLER_3_153 VPWR VGND sg13g2_fill_1
Xhold4 _0331_ VPWR VGND net410 sg13g2_dlygate4sd3_1
XFILLER_48_853 VPWR VGND sg13g2_decap_8
X_3990_ _0965_ mydesign.pe_inputs\[55\] _0914_ VPWR VGND sg13g2_nand2b_1
XFILLER_16_783 VPWR VGND sg13g2_decap_4
X_5660_ VGND VPWR net519 mydesign.pe_weights\[19\] _2448_ _2446_ sg13g2_a21oi_1
X_4611_ _0393_ _1515_ _1516_ _1517_ VPWR VGND sg13g2_nor3_2
XFILLER_30_241 VPWR VGND sg13g2_fill_2
X_5591_ _2382_ _2373_ _2383_ VPWR VGND sg13g2_xor2_1
X_4542_ _1452_ _1440_ _1453_ VPWR VGND sg13g2_xor2_1
X_6097__300 VPWR VGND net300 sg13g2_tiehi
XFILLER_7_492 VPWR VGND sg13g2_fill_1
Xhold426 mydesign.accum\[3\] VPWR VGND net1045 sg13g2_dlygate4sd3_1
Xhold415 _0200_ VPWR VGND net1034 sg13g2_dlygate4sd3_1
X_4473_ _1396_ net977 _1382_ VPWR VGND sg13g2_xnor2_1
Xhold404 _0228_ VPWR VGND net1023 sg13g2_dlygate4sd3_1
Xhold448 mydesign.pe_weights\[51\] VPWR VGND net1067 sg13g2_dlygate4sd3_1
X_3424_ VGND VPWR _0466_ _0467_ _0073_ _0468_ sg13g2_a21oi_1
Xhold459 net11 VPWR VGND net1078 sg13g2_dlygate4sd3_1
Xhold437 _0319_ VPWR VGND net1056 sg13g2_dlygate4sd3_1
X_6143_ net208 VGND VPWR _0369_ mydesign.weights\[0\]\[13\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3355_ net834 net755 _0405_ VPWR VGND sg13g2_nor2b_2
X_3286_ net614 VPWR _2686_ VGND _2620_ _2657_ sg13g2_o21ai_1
X_6074_ net136 VGND VPWR net759 mydesign.accum\[16\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_5025_ _1877_ _1875_ _1874_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_886 VPWR VGND sg13g2_decap_8
XFILLER_0_1020 VPWR VGND sg13g2_decap_8
XFILLER_26_558 VPWR VGND sg13g2_decap_8
XFILLER_13_208 VPWR VGND sg13g2_fill_2
XFILLER_34_580 VPWR VGND sg13g2_decap_8
X_5927_ net303 VGND VPWR _0153_ mydesign.pe_weights\[45\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_6067__192 VPWR VGND net192 sg13g2_tiehi
X_5858_ net57 VGND VPWR net809 mydesign.pe_weights\[60\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
X_4809_ net533 net529 mydesign.accum\[51\] _1688_ VPWR VGND sg13g2_nand3_1
X_5789_ net161 VGND VPWR net668 mydesign.inputs\[2\]\[10\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_48_149 VPWR VGND sg13g2_decap_4
XFILLER_28_30 VPWR VGND sg13g2_fill_2
XFILLER_28_41 VPWR VGND sg13g2_fill_2
XFILLER_28_52 VPWR VGND sg13g2_fill_2
XFILLER_45_856 VPWR VGND sg13g2_decap_8
XFILLER_8_234 VPWR VGND sg13g2_fill_1
XFILLER_9_768 VPWR VGND sg13g2_fill_2
XFILLER_4_440 VPWR VGND sg13g2_decap_4
X_3140_ VPWR _2581_ net1027 VGND sg13g2_inv_1
XFILLER_48_650 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_fill_2
XFILLER_36_801 VPWR VGND sg13g2_fill_2
XFILLER_35_311 VPWR VGND sg13g2_fill_2
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
XFILLER_35_333 VPWR VGND sg13g2_fill_2
XFILLER_35_388 VPWR VGND sg13g2_decap_8
X_3973_ _0949_ mydesign.pe_inputs\[54\] _0914_ VPWR VGND sg13g2_nand2b_1
X_5712_ net802 _2485_ _2481_ _0344_ VPWR VGND sg13g2_mux2_1
X_5643_ _2411_ mydesign.accum\[5\] _2432_ VPWR VGND sg13g2_xor2_1
X_6060__218 VPWR VGND net218 sg13g2_tiehi
X_5574_ _2364_ _2366_ _2367_ VPWR VGND sg13g2_nor2_1
X_6140__264 VPWR VGND net264 sg13g2_tiehi
Xhold201 mydesign.weights\[3\]\[11\] VPWR VGND net820 sg13g2_dlygate4sd3_1
X_4525_ net464 VPWR _1437_ VGND net566 net873 sg13g2_o21ai_1
Xhold234 mydesign.weights\[3\]\[10\] VPWR VGND net853 sg13g2_dlygate4sd3_1
Xhold223 mydesign.load_counter\[0\] VPWR VGND net842 sg13g2_dlygate4sd3_1
Xhold212 _0258_ VPWR VGND net831 sg13g2_dlygate4sd3_1
Xhold278 _0157_ VPWR VGND net897 sg13g2_dlygate4sd3_1
Xhold245 mydesign.accum\[35\] VPWR VGND net864 sg13g2_dlygate4sd3_1
Xhold256 mydesign.accum\[73\] VPWR VGND net875 sg13g2_dlygate4sd3_1
Xhold267 mydesign.accum\[76\] VPWR VGND net886 sg13g2_dlygate4sd3_1
X_4456_ _1380_ VPWR _1381_ VGND net583 net905 sg13g2_o21ai_1
Xhold289 _0205_ VPWR VGND net908 sg13g2_dlygate4sd3_1
X_4387_ _1315_ _1298_ _1314_ VPWR VGND sg13g2_nand2_1
X_3407_ net515 mydesign.accum\[116\] mydesign.accum\[84\] mydesign.accum\[52\] mydesign.accum\[20\]
+ net508 _0453_ VPWR VGND sg13g2_mux4_1
X_3338_ net541 net546 _0392_ VPWR VGND sg13g2_nor2b_2
X_6126_ net24 VGND VPWR net724 mydesign.weights\[0\]\[24\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3269_ VGND VPWR _2517_ _2673_ _0032_ _2677_ sg13g2_a21oi_1
XFILLER_22_1010 VPWR VGND sg13g2_decap_8
X_6057_ net230 VGND VPWR _0283_ mydesign.pe_inputs\[15\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_5008_ _1859_ _1858_ _1861_ VPWR VGND sg13g2_xor2_1
XFILLER_38_193 VPWR VGND sg13g2_fill_2
XFILLER_30_31 VPWR VGND sg13g2_fill_2
XFILLER_2_999 VPWR VGND sg13g2_decap_8
XFILLER_49_447 VPWR VGND sg13g2_decap_8
XFILLER_39_84 VPWR VGND sg13g2_fill_1
XFILLER_39_73 VPWR VGND sg13g2_fill_1
X_5876__397 VPWR VGND net397 sg13g2_tiehi
XFILLER_18_823 VPWR VGND sg13g2_decap_4
XFILLER_36_119 VPWR VGND sg13g2_fill_2
XFILLER_45_653 VPWR VGND sg13g2_decap_8
XFILLER_29_182 VPWR VGND sg13g2_decap_8
X_6128__384 VPWR VGND net384 sg13g2_tiehi
XFILLER_41_881 VPWR VGND sg13g2_decap_8
X_4310_ _1251_ mydesign.accum\[85\] net539 mydesign.pe_inputs\[46\] VPWR VGND sg13g2_and3_1
X_5290_ _2118_ _2102_ _2116_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_1010 VPWR VGND sg13g2_decap_8
X_4241_ _1186_ mydesign.pe_weights\[56\] mydesign.pe_inputs\[45\] VPWR VGND sg13g2_nand2_1
X_4172_ _1129_ _1121_ _1130_ VPWR VGND sg13g2_xor2_1
X_3123_ VPWR _2564_ net539 VGND sg13g2_inv_1
XFILLER_48_491 VPWR VGND sg13g2_fill_2
XFILLER_24_804 VPWR VGND sg13g2_fill_2
X_3956_ VGND VPWR _2553_ net486 _0139_ _0934_ sg13g2_a21oi_1
X_5626_ _2416_ _2413_ _2414_ VPWR VGND sg13g2_xnor2_1
X_3887_ VGND VPWR _0855_ _0872_ _0876_ _0871_ sg13g2_a21oi_1
X_5557_ _2355_ net606 _2354_ VPWR VGND sg13g2_nand2_2
X_4508_ _1419_ _1418_ _1421_ VPWR VGND sg13g2_xor2_1
X_5488_ _2276_ _2290_ _2291_ VPWR VGND sg13g2_and2_1
X_4439_ _1364_ mydesign.pe_weights\[54\] mydesign.pe_inputs\[43\] VPWR VGND sg13g2_nand2_1
Xfanout500 _2516_ net500 VPWR VGND sg13g2_buf_8
Xfanout533 net789 net533 VPWR VGND sg13g2_buf_8
Xfanout511 net518 net511 VPWR VGND sg13g2_buf_8
Xfanout522 net1098 net522 VPWR VGND sg13g2_buf_8
Xfanout544 net545 net544 VPWR VGND sg13g2_buf_8
Xfanout566 net571 net566 VPWR VGND sg13g2_buf_8
Xfanout555 net556 net555 VPWR VGND sg13g2_buf_1
XFILLER_47_929 VPWR VGND sg13g2_decap_8
Xfanout588 net589 net588 VPWR VGND sg13g2_buf_8
Xfanout599 _2629_ net599 VPWR VGND sg13g2_buf_8
Xfanout577 net578 net577 VPWR VGND sg13g2_buf_8
X_6109_ net216 VGND VPWR _0335_ mydesign.weights\[1\]\[19\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_6112__196 VPWR VGND net196 sg13g2_tiehi
XFILLER_15_848 VPWR VGND sg13g2_fill_1
XFILLER_25_31 VPWR VGND sg13g2_fill_1
XFILLER_30_829 VPWR VGND sg13g2_fill_1
XFILLER_22_391 VPWR VGND sg13g2_decap_8
XFILLER_6_513 VPWR VGND sg13g2_fill_2
XFILLER_10_575 VPWR VGND sg13g2_decap_4
XFILLER_41_85 VPWR VGND sg13g2_fill_2
XFILLER_6_546 VPWR VGND sg13g2_fill_2
XFILLER_2_730 VPWR VGND sg13g2_fill_2
XFILLER_2_763 VPWR VGND sg13g2_fill_1
XFILLER_1_251 VPWR VGND sg13g2_fill_2
XFILLER_37_9 VPWR VGND sg13g2_fill_1
XFILLER_49_200 VPWR VGND sg13g2_fill_2
XFILLER_37_439 VPWR VGND sg13g2_decap_8
X_3810_ net630 VPWR _0805_ VGND net491 _0804_ sg13g2_o21ai_1
X_4790_ mydesign.pe_weights\[42\] net529 mydesign.accum\[50\] _1670_ VPWR VGND sg13g2_nand3_1
X_3741_ _0749_ _0748_ _0747_ VPWR VGND sg13g2_nand2b_1
XFILLER_9_362 VPWR VGND sg13g2_fill_1
X_3672_ _0684_ _0666_ _0682_ VPWR VGND sg13g2_xnor2_1
X_5411_ net593 VPWR _2224_ VGND _2222_ _2223_ sg13g2_o21ai_1
X_5342_ _2156_ _2153_ _2158_ VPWR VGND sg13g2_xor2_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_5_590 VPWR VGND sg13g2_fill_1
X_5273_ _2102_ _2100_ _2101_ VPWR VGND sg13g2_nand2b_1
X_4224_ net626 VPWR _1176_ VGND net981 net438 sg13g2_o21ai_1
X_4155_ _1114_ _1097_ _1112_ _1113_ VPWR VGND sg13g2_and3_1
XFILLER_46_19 VPWR VGND sg13g2_fill_2
X_3106_ _2547_ net529 VPWR VGND sg13g2_inv_2
X_4086_ _1054_ _0394_ mydesign.inputs\[1\]\[14\] net461 mydesign.inputs\[1\]\[22\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_37_973 VPWR VGND sg13g2_decap_8
XFILLER_24_678 VPWR VGND sg13g2_fill_2
XFILLER_11_339 VPWR VGND sg13g2_decap_4
X_4988_ _1833_ _1841_ _1842_ VPWR VGND sg13g2_nor2_1
X_3939_ net628 VPWR _0920_ VGND net486 _0919_ sg13g2_o21ai_1
XFILLER_20_840 VPWR VGND sg13g2_fill_2
X_5609_ _2400_ _2389_ _2399_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_11 VPWR VGND sg13g2_decap_8
X_6042__290 VPWR VGND net290 sg13g2_tiehi
X_5942__273 VPWR VGND net273 sg13g2_tiehi
XFILLER_47_726 VPWR VGND sg13g2_decap_8
XFILLER_4_1018 VPWR VGND sg13g2_decap_8
XFILLER_43_921 VPWR VGND sg13g2_decap_8
XFILLER_15_601 VPWR VGND sg13g2_decap_4
XFILLER_28_984 VPWR VGND sg13g2_decap_8
XFILLER_14_133 VPWR VGND sg13g2_fill_2
XFILLER_43_998 VPWR VGND sg13g2_decap_8
XFILLER_14_166 VPWR VGND sg13g2_decap_4
XFILLER_35_1020 VPWR VGND sg13g2_decap_8
XFILLER_7_833 VPWR VGND sg13g2_decap_8
XFILLER_42_1024 VPWR VGND sg13g2_decap_4
XFILLER_38_737 VPWR VGND sg13g2_fill_1
XFILLER_38_715 VPWR VGND sg13g2_fill_1
X_5960_ net237 VGND VPWR _0186_ mydesign.pe_weights\[38\] clknet_leaf_32_clk sg13g2_dfrbpq_2
XFILLER_18_450 VPWR VGND sg13g2_fill_2
XFILLER_19_962 VPWR VGND sg13g2_decap_8
X_5891_ net371 VGND VPWR _0117_ mydesign.pe_inputs\[53\] clknet_leaf_44_clk sg13g2_dfrbpq_2
X_4911_ net634 VPWR _1777_ VGND net526 net442 sg13g2_o21ai_1
XFILLER_34_921 VPWR VGND sg13g2_decap_8
X_5889__374 VPWR VGND net374 sg13g2_tiehi
XFILLER_21_637 VPWR VGND sg13g2_decap_8
XFILLER_33_475 VPWR VGND sg13g2_fill_2
XFILLER_34_998 VPWR VGND sg13g2_decap_8
X_4842_ _1718_ _1717_ _1720_ VPWR VGND sg13g2_xor2_1
X_4773_ VGND VPWR _2541_ net451 _0235_ _1655_ sg13g2_a21oi_1
XFILLER_21_648 VPWR VGND sg13g2_decap_4
X_3724_ mydesign.pe_inputs\[62\] _0658_ mydesign.accum\[117\] _0733_ VPWR VGND sg13g2_nand3_1
X_3655_ _0666_ _0667_ _0668_ VPWR VGND sg13g2_nor2_1
X_3586_ _0611_ _0589_ _0609_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_508 VPWR VGND sg13g2_fill_1
X_5325_ _2142_ mydesign.accum\[17\] net522 mydesign.pe_weights\[25\] VPWR VGND sg13g2_and3_2
X_5256_ _2086_ _2079_ _2084_ VPWR VGND sg13g2_xnor2_1
X_4207_ _1163_ _1147_ _1149_ VPWR VGND sg13g2_nand2_1
XFILLER_29_704 VPWR VGND sg13g2_decap_8
X_5187_ VGND VPWR _2525_ net494 _0283_ _2021_ sg13g2_a21oi_1
X_4138_ _1097_ _1087_ _1089_ VPWR VGND sg13g2_nand2_1
XFILLER_44_729 VPWR VGND sg13g2_decap_8
X_4069_ _1040_ _1030_ _1039_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_910 VPWR VGND sg13g2_fill_2
XFILLER_37_792 VPWR VGND sg13g2_fill_1
X_6081__60 VPWR VGND net60 sg13g2_tiehi
XFILLER_19_1004 VPWR VGND sg13g2_decap_8
XFILLER_25_987 VPWR VGND sg13g2_decap_8
XFILLER_40_924 VPWR VGND sg13g2_decap_8
XFILLER_3_335 VPWR VGND sg13g2_fill_1
XFILLER_47_512 VPWR VGND sg13g2_decap_4
XFILLER_47_567 VPWR VGND sg13g2_fill_1
XFILLER_35_729 VPWR VGND sg13g2_fill_1
XFILLER_43_795 VPWR VGND sg13g2_decap_8
XFILLER_16_998 VPWR VGND sg13g2_decap_8
XFILLER_31_957 VPWR VGND sg13g2_decap_8
XFILLER_30_478 VPWR VGND sg13g2_decap_8
XFILLER_11_681 VPWR VGND sg13g2_fill_1
X_3440_ net511 mydesign.accum\[127\] mydesign.accum\[95\] mydesign.accum\[63\] mydesign.accum\[31\]
+ net505 _0483_ VPWR VGND sg13g2_mux4_1
X_3371_ net515 mydesign.accum\[113\] mydesign.accum\[81\] mydesign.accum\[49\] mydesign.accum\[17\]
+ net508 _0420_ VPWR VGND sg13g2_mux4_1
X_5110_ _1951_ _1942_ _1952_ VPWR VGND sg13g2_xor2_1
X_6090_ net360 VGND VPWR _0316_ mydesign.accum\[12\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_6056__234 VPWR VGND net234 sg13g2_tiehi
X_5041_ VGND VPWR _2532_ net443 _0268_ _1890_ sg13g2_a21oi_1
XFILLER_25_206 VPWR VGND sg13g2_fill_2
XFILLER_19_792 VPWR VGND sg13g2_fill_2
X_5943_ net271 VGND VPWR _0169_ mydesign.pe_weights\[41\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_5874_ net25 VGND VPWR _0100_ mydesign.pe_weights\[56\] clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_22_924 VPWR VGND sg13g2_decap_4
XFILLER_22_968 VPWR VGND sg13g2_decap_8
X_4825_ VGND VPWR net582 _1702_ _0239_ _1703_ sg13g2_a21oi_1
X_4756_ net470 VPWR _1647_ VGND net567 net941 sg13g2_o21ai_1
XFILLER_30_990 VPWR VGND sg13g2_decap_8
X_4687_ _1557_ _1581_ _1582_ VPWR VGND sg13g2_nor2b_1
X_3707_ _0715_ _0713_ _0717_ VPWR VGND sg13g2_xor2_1
X_3638_ net630 VPWR _0654_ VGND net487 _0653_ sg13g2_o21ai_1
X_3569_ _0575_ _0572_ _0593_ _0595_ VPWR VGND sg13g2_a21o_1
XFILLER_1_817 VPWR VGND sg13g2_fill_1
X_5308_ _2133_ net660 _2131_ VPWR VGND sg13g2_nand2_1
X_6035__318 VPWR VGND net318 sg13g2_tiehi
X_5239_ _2067_ _2068_ _2052_ _2070_ VPWR VGND sg13g2_nand3_1
XFILLER_29_512 VPWR VGND sg13g2_fill_2
XFILLER_44_504 VPWR VGND sg13g2_fill_1
XFILLER_24_283 VPWR VGND sg13g2_fill_2
XFILLER_12_478 VPWR VGND sg13g2_fill_1
XFILLER_4_666 VPWR VGND sg13g2_decap_4
XFILLER_4_699 VPWR VGND sg13g2_fill_2
XFILLER_4_688 VPWR VGND sg13g2_decap_8
XFILLER_48_832 VPWR VGND sg13g2_decap_8
Xhold5 mydesign.weights\[3\]\[4\] VPWR VGND net411 sg13g2_dlygate4sd3_1
XFILLER_0_894 VPWR VGND sg13g2_decap_8
XFILLER_16_740 VPWR VGND sg13g2_decap_8
X_5886__377 VPWR VGND net377 sg13g2_tiehi
X_4610_ mydesign.inputs\[2\]\[12\] net550 _1516_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_787 VPWR VGND sg13g2_decap_4
X_5590_ _2382_ _2374_ _2380_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_297 VPWR VGND sg13g2_decap_8
X_4541_ _1452_ _1428_ _1450_ VPWR VGND sg13g2_xnor2_1
Xhold416 mydesign.accum\[21\] VPWR VGND net1035 sg13g2_dlygate4sd3_1
XFILLER_8_994 VPWR VGND sg13g2_decap_8
Xhold405 mydesign.pe_inputs\[53\] VPWR VGND net1024 sg13g2_dlygate4sd3_1
X_4472_ VGND VPWR _1371_ _1386_ _1395_ _1385_ sg13g2_a21oi_1
Xhold427 mydesign.pe_inputs\[59\] VPWR VGND net1046 sg13g2_dlygate4sd3_1
Xhold449 mydesign.accum\[4\] VPWR VGND net1068 sg13g2_dlygate4sd3_1
Xhold438 mydesign.accum\[1\] VPWR VGND net1057 sg13g2_dlygate4sd3_1
X_3423_ net622 VPWR _0468_ VGND net1080 net431 sg13g2_o21ai_1
X_6142_ net232 VGND VPWR _0368_ mydesign.weights\[0\]\[12\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3354_ net513 mydesign.accum\[96\] mydesign.accum\[64\] mydesign.accum\[32\] mydesign.accum\[0\]
+ net506 _0404_ VPWR VGND sg13g2_mux4_1
XFILLER_31_0 VPWR VGND sg13g2_fill_1
X_3285_ _2670_ net778 _2685_ _0040_ VPWR VGND sg13g2_mux2_1
X_6073_ net144 VGND VPWR net1001 mydesign.pe_inputs\[11\] clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_39_843 VPWR VGND sg13g2_fill_1
XFILLER_39_832 VPWR VGND sg13g2_fill_1
X_5024_ _1875_ _1874_ _1876_ VPWR VGND sg13g2_nor2b_1
X_5926_ net305 VGND VPWR _0152_ mydesign.pe_weights\[44\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_5857_ net59 VGND VPWR _0083_ mydesign.pe_inputs\[63\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_4808_ _1687_ mydesign.pe_weights\[42\] mydesign.pe_inputs\[29\] VPWR VGND sg13g2_nand2_1
XFILLER_6_909 VPWR VGND sg13g2_fill_2
XFILLER_10_949 VPWR VGND sg13g2_decap_8
XFILLER_22_798 VPWR VGND sg13g2_decap_8
X_5788_ net162 VGND VPWR net421 mydesign.inputs\[2\]\[9\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_5_419 VPWR VGND sg13g2_fill_2
X_4739_ VGND VPWR net535 _1537_ _1631_ mydesign.accum\[62\] sg13g2_a21oi_1
XFILLER_49_629 VPWR VGND sg13g2_decap_8
XFILLER_48_117 VPWR VGND sg13g2_fill_1
XFILLER_29_353 VPWR VGND sg13g2_fill_2
XFILLER_45_835 VPWR VGND sg13g2_decap_8
X_5831__107 VPWR VGND net107 sg13g2_tiehi
XFILLER_29_386 VPWR VGND sg13g2_fill_1
XFILLER_32_518 VPWR VGND sg13g2_decap_8
XFILLER_40_540 VPWR VGND sg13g2_decap_4
XFILLER_8_202 VPWR VGND sg13g2_fill_1
XFILLER_5_986 VPWR VGND sg13g2_decap_8
XFILLER_4_485 VPWR VGND sg13g2_fill_1
XFILLER_4_474 VPWR VGND sg13g2_decap_8
XFILLER_39_128 VPWR VGND sg13g2_decap_8
XFILLER_35_345 VPWR VGND sg13g2_fill_1
XFILLER_23_518 VPWR VGND sg13g2_fill_1
XFILLER_44_890 VPWR VGND sg13g2_decap_8
X_3972_ VGND VPWR net564 _0947_ _0141_ _0948_ sg13g2_a21oi_1
X_5711_ _2520_ _2484_ _2485_ VPWR VGND sg13g2_nor2_2
X_5642_ mydesign.accum\[4\] net519 mydesign.accum\[5\] _2431_ VPWR VGND mydesign.pe_weights\[17\]
+ sg13g2_nand4_1
X_5573_ VGND VPWR mydesign.pe_inputs\[5\] net524 _2366_ mydesign.accum\[1\] sg13g2_a21oi_1
X_4524_ _1436_ _1420_ _1435_ VPWR VGND sg13g2_xnor2_1
Xhold202 _1776_ VPWR VGND net821 sg13g2_dlygate4sd3_1
X_5782__172 VPWR VGND net172 sg13g2_tiehi
Xhold235 _1774_ VPWR VGND net854 sg13g2_dlygate4sd3_1
Xhold224 mydesign.accum\[71\] VPWR VGND net843 sg13g2_dlygate4sd3_1
Xhold213 mydesign.pe_inputs\[10\] VPWR VGND net832 sg13g2_dlygate4sd3_1
Xhold246 mydesign.accum\[87\] VPWR VGND net865 sg13g2_dlygate4sd3_1
Xhold257 _0189_ VPWR VGND net876 sg13g2_dlygate4sd3_1
X_4455_ net576 VPWR _1380_ VGND _1378_ _1379_ sg13g2_o21ai_1
Xhold268 mydesign.pe_inputs\[31\] VPWR VGND net887 sg13g2_dlygate4sd3_1
Xhold279 mydesign.accum\[118\] VPWR VGND net898 sg13g2_dlygate4sd3_1
X_4386_ _1312_ _1309_ _1314_ VPWR VGND sg13g2_xor2_1
X_3406_ net518 mydesign.accum\[124\] mydesign.accum\[92\] mydesign.accum\[60\] mydesign.accum\[28\]
+ net505 _0452_ VPWR VGND sg13g2_mux4_1
X_3337_ net607 _0391_ _0063_ VPWR VGND sg13g2_nor2_1
X_6125_ net32 VGND VPWR _0351_ mydesign.weights\[1\]\[15\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_3268_ net617 VPWR _2677_ VGND net885 _2673_ sg13g2_o21ai_1
XFILLER_27_802 VPWR VGND sg13g2_fill_2
X_6056_ net234 VGND VPWR _0282_ mydesign.pe_inputs\[14\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_5007_ _1860_ _1858_ _1859_ VPWR VGND sg13g2_nand2_1
X_3199_ _2630_ VPWR _0008_ VGND _2623_ net598 sg13g2_o21ai_1
XFILLER_38_161 VPWR VGND sg13g2_fill_2
XFILLER_42_805 VPWR VGND sg13g2_decap_4
XFILLER_26_323 VPWR VGND sg13g2_fill_1
XFILLER_42_816 VPWR VGND sg13g2_fill_2
XFILLER_42_849 VPWR VGND sg13g2_decap_8
X_5909_ net338 VGND VPWR _0135_ mydesign.inputs\[0\]\[23\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_10_779 VPWR VGND sg13g2_fill_2
XFILLER_5_205 VPWR VGND sg13g2_fill_1
XFILLER_2_923 VPWR VGND sg13g2_fill_1
XFILLER_49_404 VPWR VGND sg13g2_decap_4
XFILLER_7_1016 VPWR VGND sg13g2_decap_8
XFILLER_2_978 VPWR VGND sg13g2_decap_8
XFILLER_7_1027 VPWR VGND sg13g2_fill_2
X_5952__253 VPWR VGND net253 sg13g2_tiehi
X_5853__66 VPWR VGND net66 sg13g2_tiehi
XFILLER_45_632 VPWR VGND sg13g2_decap_8
XFILLER_44_142 VPWR VGND sg13g2_fill_2
XFILLER_44_186 VPWR VGND sg13g2_fill_2
X_6015__30 VPWR VGND net30 sg13g2_tiehi
X_6087__388 VPWR VGND net388 sg13g2_tiehi
XFILLER_41_860 VPWR VGND sg13g2_decap_8
XFILLER_9_522 VPWR VGND sg13g2_fill_2
X_4240_ VGND VPWR mydesign.pe_weights\[57\] net536 _1185_ mydesign.accum\[81\] sg13g2_a21oi_1
XFILLER_5_794 VPWR VGND sg13g2_fill_2
X_4171_ _1129_ _1122_ _1127_ VPWR VGND sg13g2_xnor2_1
X_3122_ VPWR _2563_ net534 VGND sg13g2_inv_1
XFILLER_49_993 VPWR VGND sg13g2_decap_8
XFILLER_36_676 VPWR VGND sg13g2_fill_1
XFILLER_24_849 VPWR VGND sg13g2_fill_2
XFILLER_36_698 VPWR VGND sg13g2_decap_4
X_3955_ net628 VPWR _0934_ VGND net486 net428 sg13g2_o21ai_1
X_5625_ VPWR _2415_ _2414_ VGND sg13g2_inv_1
X_3886_ VGND VPWR net501 _2579_ _0128_ _0875_ sg13g2_a21oi_1
X_5929__299 VPWR VGND net299 sg13g2_tiehi
XFILLER_3_709 VPWR VGND sg13g2_decap_8
X_5556_ _2607_ _2683_ _2354_ VPWR VGND sg13g2_nor2_2
XFILLER_2_208 VPWR VGND sg13g2_fill_2
X_4507_ mydesign.pe_weights\[48\] mydesign.pe_inputs\[36\] net690 _1420_ VPWR VGND
+ _1418_ sg13g2_nand4_1
X_5487_ _2289_ _2277_ _2290_ VPWR VGND sg13g2_xor2_1
X_4438_ _1362_ _1363_ _0192_ VPWR VGND sg13g2_nor2_1
Xfanout501 net503 net501 VPWR VGND sg13g2_buf_8
Xfanout523 net524 net523 VPWR VGND sg13g2_buf_2
Xfanout512 net518 net512 VPWR VGND sg13g2_buf_8
X_4369_ _1298_ mydesign.accum\[73\] mydesign.pe_weights\[53\] net534 VPWR VGND sg13g2_and3_2
Xfanout534 net1050 net534 VPWR VGND sg13g2_buf_8
Xfanout545 net546 net545 VPWR VGND sg13g2_buf_8
Xfanout556 net557 net556 VPWR VGND sg13g2_buf_8
XFILLER_47_908 VPWR VGND sg13g2_decap_8
Xfanout567 net569 net567 VPWR VGND sg13g2_buf_8
Xfanout589 net594 net589 VPWR VGND sg13g2_buf_2
Xfanout578 net581 net578 VPWR VGND sg13g2_buf_2
X_6108_ net220 VGND VPWR _0334_ mydesign.weights\[1\]\[18\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_6039_ net302 VGND VPWR _0265_ mydesign.accum\[45\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_5835__99 VPWR VGND net99 sg13g2_tiehi
X_5850__69 VPWR VGND net69 sg13g2_tiehi
XFILLER_41_123 VPWR VGND sg13g2_decap_8
XFILLER_25_98 VPWR VGND sg13g2_fill_1
X_5908__339 VPWR VGND net339 sg13g2_tiehi
XFILLER_10_554 VPWR VGND sg13g2_fill_2
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_775 VPWR VGND sg13g2_fill_1
XFILLER_2_797 VPWR VGND sg13g2_decap_8
XFILLER_49_234 VPWR VGND sg13g2_fill_1
XFILLER_49_289 VPWR VGND sg13g2_decap_8
XFILLER_46_985 VPWR VGND sg13g2_decap_8
X_3740_ mydesign.pe_inputs\[63\] _0658_ mydesign.accum\[118\] _0748_ VPWR VGND sg13g2_nand3_1
XFILLER_20_318 VPWR VGND sg13g2_fill_2
X_3671_ _0683_ _0666_ _0682_ VPWR VGND sg13g2_nand2_1
X_5410_ VGND VPWR _2202_ _2205_ _2223_ _2221_ sg13g2_a21oi_1
X_5341_ _2153_ _2156_ _2157_ VPWR VGND sg13g2_nor2_1
X_6098__292 VPWR VGND net292 sg13g2_tiehi
X_5272_ VGND VPWR mydesign.accum\[28\] _2081_ _2101_ _2083_ sg13g2_a21oi_1
X_4223_ VGND VPWR _2570_ net438 _0165_ _1175_ sg13g2_a21oi_1
X_4154_ _1111_ _1110_ _1099_ _1113_ VPWR VGND sg13g2_a21o_1
X_4085_ _1053_ mydesign.inputs\[1\]\[18\] net496 VPWR VGND sg13g2_nand2_1
XFILLER_28_407 VPWR VGND sg13g2_decap_8
XFILLER_28_429 VPWR VGND sg13g2_fill_2
X_3105_ VPWR _2546_ net879 VGND sg13g2_inv_1
XFILLER_49_790 VPWR VGND sg13g2_decap_8
XFILLER_37_952 VPWR VGND sg13g2_decap_8
XFILLER_24_657 VPWR VGND sg13g2_decap_8
X_4987_ _1841_ _1834_ _1839_ VPWR VGND sg13g2_xnor2_1
X_3938_ _0918_ VPWR _0919_ VGND _0916_ _0917_ sg13g2_o21ai_1
X_3869_ _0859_ mydesign.pe_inputs\[58\] _0796_ VPWR VGND sg13g2_nand2_1
X_5608_ _2396_ _2390_ _2399_ VPWR VGND sg13g2_xor2_1
X_5539_ _2322_ _2338_ _2321_ _2339_ VPWR VGND sg13g2_nand3_1
XFILLER_3_539 VPWR VGND sg13g2_fill_1
XFILLER_47_705 VPWR VGND sg13g2_decap_8
XFILLER_43_900 VPWR VGND sg13g2_decap_8
XFILLER_28_963 VPWR VGND sg13g2_decap_8
XFILLER_36_53 VPWR VGND sg13g2_fill_1
XFILLER_42_421 VPWR VGND sg13g2_decap_8
XFILLER_43_977 VPWR VGND sg13g2_decap_8
XFILLER_42_476 VPWR VGND sg13g2_decap_4
XFILLER_10_340 VPWR VGND sg13g2_fill_2
XFILLER_7_856 VPWR VGND sg13g2_fill_1
XFILLER_6_377 VPWR VGND sg13g2_decap_8
XFILLER_6_388 VPWR VGND sg13g2_fill_2
X_5804__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_42_1003 VPWR VGND sg13g2_decap_8
X_6132__348 VPWR VGND net348 sg13g2_tiehi
XFILLER_19_941 VPWR VGND sg13g2_decap_8
XFILLER_18_462 VPWR VGND sg13g2_fill_1
XFILLER_34_900 VPWR VGND sg13g2_decap_8
XFILLER_46_782 VPWR VGND sg13g2_decap_8
X_4910_ VGND VPWR _1767_ _1775_ _0251_ net821 sg13g2_a21oi_1
X_5890_ net373 VGND VPWR _0116_ mydesign.pe_inputs\[52\] clknet_leaf_44_clk sg13g2_dfrbpq_2
XFILLER_34_977 VPWR VGND sg13g2_decap_8
X_4841_ _1719_ _1717_ _1718_ VPWR VGND sg13g2_nand2_1
XFILLER_20_137 VPWR VGND sg13g2_decap_8
X_4772_ net638 VPWR _1655_ VGND net527 net451 sg13g2_o21ai_1
X_3723_ _0732_ mydesign.pe_inputs\[63\] _0653_ VPWR VGND sg13g2_nand2_1
X_3654_ _0667_ _0663_ _0665_ _0643_ mydesign.pe_inputs\[61\] VPWR VGND sg13g2_a22oi_1
X_3585_ _0589_ _0609_ _0610_ VPWR VGND sg13g2_nor2_1
X_5324_ VGND VPWR net758 _2140_ _0300_ _2141_ sg13g2_a21oi_1
X_5255_ _2085_ _2079_ _2084_ VPWR VGND sg13g2_nand2_1
X_4206_ _1149_ _1160_ _1162_ VPWR VGND sg13g2_nor2_1
X_5186_ net625 VPWR _2021_ VGND net487 _2020_ sg13g2_o21ai_1
X_4137_ VGND VPWR _1076_ _1092_ _1096_ _1091_ sg13g2_a21oi_1
XFILLER_44_708 VPWR VGND sg13g2_decap_8
X_4068_ _1039_ net940 _1038_ VPWR VGND sg13g2_xnor2_1
XFILLER_40_903 VPWR VGND sg13g2_decap_8
XFILLER_24_443 VPWR VGND sg13g2_decap_8
XFILLER_25_966 VPWR VGND sg13g2_decap_8
XFILLER_20_682 VPWR VGND sg13g2_fill_2
XFILLER_22_44 VPWR VGND sg13g2_fill_1
XFILLER_4_859 VPWR VGND sg13g2_fill_2
XFILLER_3_358 VPWR VGND sg13g2_decap_4
XFILLER_26_1009 VPWR VGND sg13g2_decap_8
XFILLER_16_977 VPWR VGND sg13g2_decap_8
XFILLER_43_774 VPWR VGND sg13g2_decap_8
XFILLER_30_413 VPWR VGND sg13g2_decap_4
XFILLER_31_936 VPWR VGND sg13g2_decap_8
XFILLER_10_170 VPWR VGND sg13g2_fill_1
X_3370_ VGND VPWR net458 _0418_ _0419_ _2698_ sg13g2_a21oi_1
XFILLER_2_380 VPWR VGND sg13g2_decap_8
X_5040_ net634 VPWR _1890_ VGND net903 net443 sg13g2_o21ai_1
XFILLER_25_218 VPWR VGND sg13g2_fill_1
X_5942_ net273 VGND VPWR _0168_ mydesign.pe_weights\[40\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_6063__206 VPWR VGND net206 sg13g2_tiehi
XFILLER_22_914 VPWR VGND sg13g2_decap_4
X_5873_ net27 VGND VPWR _0099_ mydesign.pe_inputs\[59\] clknet_leaf_7_clk sg13g2_dfrbpq_2
XFILLER_34_785 VPWR VGND sg13g2_decap_8
XFILLER_22_947 VPWR VGND sg13g2_decap_8
X_4824_ net479 VPWR _1703_ VGND net582 net969 sg13g2_o21ai_1
X_4755_ _1646_ _1642_ _1645_ VPWR VGND sg13g2_xnor2_1
X_3706_ _0713_ _0715_ _0716_ VPWR VGND sg13g2_nor2_1
X_4686_ _1581_ _1576_ _1580_ VPWR VGND sg13g2_xnor2_1
X_3637_ _0650_ VPWR _0653_ VGND net542 _0652_ sg13g2_o21ai_1
X_3568_ _0575_ _0593_ _0572_ _0594_ VPWR VGND sg13g2_nand3_1
XFILLER_0_317 VPWR VGND sg13g2_decap_8
XFILLER_1_829 VPWR VGND sg13g2_decap_8
X_5307_ _2132_ VPWR _0292_ VGND net603 _2130_ sg13g2_o21ai_1
X_3499_ net467 VPWR _0529_ VGND net721 _0528_ sg13g2_o21ai_1
X_5238_ _2069_ _2067_ _2068_ VPWR VGND sg13g2_nand2_1
X_5169_ _2006_ mydesign.inputs\[3\]\[9\] net549 VPWR VGND sg13g2_nand2b_1
X_5911__335 VPWR VGND net335 sg13g2_tiehi
XFILLER_12_413 VPWR VGND sg13g2_decap_8
XFILLER_33_21 VPWR VGND sg13g2_fill_2
XFILLER_33_43 VPWR VGND sg13g2_decap_4
XFILLER_8_406 VPWR VGND sg13g2_decap_4
XFILLER_32_1013 VPWR VGND sg13g2_decap_8
XFILLER_48_811 VPWR VGND sg13g2_decap_8
XFILLER_0_873 VPWR VGND sg13g2_decap_8
Xhold6 _0112_ VPWR VGND net412 sg13g2_dlygate4sd3_1
XFILLER_48_888 VPWR VGND sg13g2_decap_8
XFILLER_47_332 VPWR VGND sg13g2_decap_4
XFILLER_35_505 VPWR VGND sg13g2_decap_8
XFILLER_30_243 VPWR VGND sg13g2_fill_1
X_5962__233 VPWR VGND net233 sg13g2_tiehi
XFILLER_12_991 VPWR VGND sg13g2_decap_8
XFILLER_8_973 VPWR VGND sg13g2_decap_8
XFILLER_8_951 VPWR VGND sg13g2_fill_2
X_4540_ _1451_ _1428_ _1450_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_10_clk clknet_3_0__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
Xhold417 mydesign.pe_inputs\[54\] VPWR VGND net1036 sg13g2_dlygate4sd3_1
Xhold406 mydesign.pe_weights\[23\] VPWR VGND net1025 sg13g2_dlygate4sd3_1
X_4471_ _1391_ VPWR _1394_ VGND _1374_ _1387_ sg13g2_o21ai_1
Xhold439 _0325_ VPWR VGND net1058 sg13g2_dlygate4sd3_1
Xhold428 _0119_ VPWR VGND net1047 sg13g2_dlygate4sd3_1
X_3422_ VGND VPWR net457 _0465_ _0467_ _0462_ sg13g2_a21oi_1
X_6141_ net248 VGND VPWR net871 mydesign.weights\[3\]\[15\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3353_ mydesign.out\[0\] mydesign.out\[1\] _0403_ VPWR VGND sg13g2_and2_1
X_3284_ _2669_ net776 _2685_ _0039_ VPWR VGND sg13g2_mux2_1
X_6072_ net168 VGND VPWR _0298_ mydesign.pe_inputs\[10\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_5023_ _1855_ VPWR _1875_ VGND _1854_ _1857_ sg13g2_o21ai_1
X_5925_ net307 VGND VPWR _0151_ mydesign.pe_inputs\[47\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_5856_ net61 VGND VPWR _0082_ mydesign.pe_inputs\[62\] clknet_leaf_20_clk sg13g2_dfrbpq_2
XFILLER_16_1019 VPWR VGND sg13g2_decap_8
XFILLER_22_766 VPWR VGND sg13g2_fill_2
X_4807_ _1686_ mydesign.pe_weights\[41\] mydesign.pe_inputs\[30\] VPWR VGND sg13g2_nand2_1
XFILLER_21_265 VPWR VGND sg13g2_decap_4
X_5787_ net163 VGND VPWR net424 mydesign.inputs\[2\]\[8\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_4738_ _1626_ VPWR _1630_ VGND _1613_ _1627_ sg13g2_o21ai_1
X_4669_ _1565_ _1555_ _1563_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_608 VPWR VGND sg13g2_decap_8
X_5939__279 VPWR VGND net279 sg13g2_tiehi
XFILLER_28_54 VPWR VGND sg13g2_fill_1
XFILLER_45_814 VPWR VGND sg13g2_decap_8
XFILLER_17_527 VPWR VGND sg13g2_decap_4
XFILLER_44_324 VPWR VGND sg13g2_fill_1
XFILLER_44_75 VPWR VGND sg13g2_decap_8
XFILLER_40_530 VPWR VGND sg13g2_fill_1
XFILLER_9_704 VPWR VGND sg13g2_decap_8
XFILLER_5_921 VPWR VGND sg13g2_fill_1
XFILLER_5_965 VPWR VGND sg13g2_decap_8
XFILLER_10_6 VPWR VGND sg13g2_fill_1
XFILLER_48_685 VPWR VGND sg13g2_decap_8
XFILLER_35_313 VPWR VGND sg13g2_fill_1
XFILLER_36_836 VPWR VGND sg13g2_fill_2
XFILLER_39_1019 VPWR VGND sg13g2_decap_8
XFILLER_35_335 VPWR VGND sg13g2_fill_1
X_3971_ net464 VPWR _0948_ VGND net564 net1007 sg13g2_o21ai_1
XFILLER_35_357 VPWR VGND sg13g2_decap_4
X_5710_ net432 _2482_ _2483_ _2484_ VPWR VGND sg13g2_nor3_2
X_5641_ _2417_ VPWR _2430_ VGND _2413_ _2415_ sg13g2_o21ai_1
X_5572_ mydesign.pe_inputs\[5\] net524 mydesign.accum\[1\] _2365_ VPWR VGND sg13g2_nand3_1
X_4523_ _1435_ _1416_ _1433_ VPWR VGND sg13g2_xnor2_1
Xhold203 _0251_ VPWR VGND net822 sg13g2_dlygate4sd3_1
Xhold225 mydesign.weights\[3\]\[8\] VPWR VGND net844 sg13g2_dlygate4sd3_1
Xhold214 _0310_ VPWR VGND net833 sg13g2_dlygate4sd3_1
Xhold236 _0250_ VPWR VGND net855 sg13g2_dlygate4sd3_1
X_4454_ VGND VPWR _1358_ _1361_ _1379_ _1377_ sg13g2_a21oi_1
Xhold269 _0231_ VPWR VGND net888 sg13g2_dlygate4sd3_1
Xhold258 mydesign.accum\[114\] VPWR VGND net877 sg13g2_dlygate4sd3_1
Xhold247 mydesign.accum\[60\] VPWR VGND net866 sg13g2_dlygate4sd3_1
X_4385_ _1309_ _1312_ _1313_ VPWR VGND sg13g2_nor2_1
X_3405_ net513 mydesign.accum\[108\] mydesign.accum\[76\] mydesign.accum\[44\] mydesign.accum\[12\]
+ net508 _0451_ VPWR VGND sg13g2_mux4_1
X_3336_ _0391_ net461 _0387_ _0389_ net546 VPWR VGND sg13g2_a22oi_1
X_6124_ net40 VGND VPWR _0350_ mydesign.weights\[1\]\[14\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_6055_ net238 VGND VPWR _0281_ mydesign.pe_inputs\[13\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_5847__75 VPWR VGND net75 sg13g2_tiehi
X_3267_ VGND VPWR _2518_ _2673_ _0031_ _2676_ sg13g2_a21oi_1
X_5006_ _1836_ VPWR _1859_ VGND _1835_ _1838_ sg13g2_o21ai_1
X_3198_ _2631_ net4 net620 VPWR VGND sg13g2_nand2_2
XFILLER_27_869 VPWR VGND sg13g2_fill_2
XFILLER_42_828 VPWR VGND sg13g2_decap_8
XFILLER_35_880 VPWR VGND sg13g2_decap_8
X_5908_ net339 VGND VPWR _0134_ mydesign.inputs\[0\]\[22\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5839_ net91 VGND VPWR _0065_ mydesign.cp2\[0\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_10_747 VPWR VGND sg13g2_fill_2
XFILLER_2_957 VPWR VGND sg13g2_decap_8
XFILLER_39_20 VPWR VGND sg13g2_decap_4
XFILLER_17_335 VPWR VGND sg13g2_decap_8
XFILLER_45_688 VPWR VGND sg13g2_decap_8
XFILLER_40_360 VPWR VGND sg13g2_decap_8
X_4170_ _1128_ _1122_ _1127_ VPWR VGND sg13g2_nand2_1
X_3121_ VPWR _2562_ net899 VGND sg13g2_inv_1
XFILLER_49_972 VPWR VGND sg13g2_decap_8
XFILLER_48_493 VPWR VGND sg13g2_fill_1
XFILLER_35_143 VPWR VGND sg13g2_decap_8
XFILLER_17_891 VPWR VGND sg13g2_fill_2
X_3954_ _0930_ _0931_ _0932_ _0933_ VPWR VGND sg13g2_or3_1
X_3885_ net465 VPWR _0875_ VGND net501 _0874_ sg13g2_o21ai_1
XFILLER_32_894 VPWR VGND sg13g2_decap_8
X_5624_ _2393_ VPWR _2414_ VGND _2391_ _2394_ sg13g2_o21ai_1
X_5555_ VGND VPWR net592 _2352_ _0319_ _2353_ sg13g2_a21oi_1
X_4506_ mydesign.pe_weights\[48\] mydesign.pe_inputs\[36\] net690 _1419_ VPWR VGND
+ sg13g2_nand3_1
X_5899__355 VPWR VGND net355 sg13g2_tiehi
X_5486_ _2289_ _2265_ _2287_ VPWR VGND sg13g2_xnor2_1
X_4437_ net474 VPWR _1363_ VGND net573 net886 sg13g2_o21ai_1
Xfanout502 net503 net502 VPWR VGND sg13g2_buf_8
Xfanout524 net903 net524 VPWR VGND sg13g2_buf_1
Xfanout513 net514 net513 VPWR VGND sg13g2_buf_8
X_4368_ VGND VPWR net684 _1296_ _0188_ _1297_ sg13g2_a21oi_1
Xfanout546 net1088 net546 VPWR VGND sg13g2_buf_8
Xfanout557 mydesign.cp\[0\] net557 VPWR VGND sg13g2_buf_8
X_6107_ net224 VGND VPWR _0333_ mydesign.weights\[1\]\[17\] clknet_leaf_11_clk sg13g2_dfrbpq_1
Xfanout535 net927 net535 VPWR VGND sg13g2_buf_8
X_4299_ _1218_ _1220_ _1239_ _1241_ VPWR VGND sg13g2_or3_1
Xfanout579 net580 net579 VPWR VGND sg13g2_buf_8
Xfanout568 net569 net568 VPWR VGND sg13g2_buf_1
X_3319_ _2620_ _2648_ _2600_ _0379_ VPWR VGND sg13g2_nand3_1
X_6038_ net306 VGND VPWR _0264_ mydesign.accum\[44\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_27_622 VPWR VGND sg13g2_fill_1
XFILLER_27_644 VPWR VGND sg13g2_decap_8
XFILLER_26_132 VPWR VGND sg13g2_fill_1
XFILLER_41_179 VPWR VGND sg13g2_decap_4
XFILLER_6_515 VPWR VGND sg13g2_fill_1
XFILLER_41_87 VPWR VGND sg13g2_fill_1
XFILLER_2_732 VPWR VGND sg13g2_fill_1
XFILLER_29_1007 VPWR VGND sg13g2_decap_8
XFILLER_49_246 VPWR VGND sg13g2_fill_1
XFILLER_38_909 VPWR VGND sg13g2_decap_8
XFILLER_46_964 VPWR VGND sg13g2_decap_8
XFILLER_45_496 VPWR VGND sg13g2_fill_2
XFILLER_14_861 VPWR VGND sg13g2_fill_1
X_3670_ _0682_ _0673_ _0680_ VPWR VGND sg13g2_xnor2_1
X_6059__222 VPWR VGND net222 sg13g2_tiehi
X_5340_ _2156_ _2154_ _2155_ VPWR VGND sg13g2_nand2_1
X_5271_ _2099_ _2096_ _2100_ VPWR VGND sg13g2_xor2_1
X_4222_ net630 VPWR _1175_ VGND net899 net438 sg13g2_o21ai_1
X_4153_ _1110_ _1111_ _1099_ _1112_ VPWR VGND sg13g2_nand3_1
XFILLER_29_909 VPWR VGND sg13g2_decap_8
X_4084_ VGND VPWR _2570_ net488 _0149_ _1052_ sg13g2_a21oi_1
X_3104_ VPWR _2545_ net887 VGND sg13g2_inv_1
XFILLER_37_931 VPWR VGND sg13g2_decap_8
XFILLER_36_441 VPWR VGND sg13g2_fill_1
X_4986_ _1834_ _1839_ _1840_ VPWR VGND sg13g2_and2_1
X_3937_ _0918_ _0395_ mydesign.weights\[3\]\[13\] net454 mydesign.weights\[3\]\[1\]
+ VPWR VGND sg13g2_a22oi_1
X_5907__340 VPWR VGND net340 sg13g2_tiehi
X_3868_ _0840_ VPWR _0858_ VGND _0838_ _0841_ sg13g2_o21ai_1
X_5607_ _2390_ _2396_ _2398_ VPWR VGND sg13g2_nor2_1
X_3799_ _0795_ _0392_ _0794_ VPWR VGND sg13g2_nand2_2
XFILLER_11_57 VPWR VGND sg13g2_fill_2
X_5538_ _2338_ _2335_ _2336_ VPWR VGND sg13g2_xnor2_1
X_6038__306 VPWR VGND net306 sg13g2_tiehi
XFILLER_2_8 VPWR VGND sg13g2_fill_2
X_5469_ _2273_ _2257_ _2272_ VPWR VGND sg13g2_xnor2_1
XFILLER_46_249 VPWR VGND sg13g2_fill_2
XFILLER_28_942 VPWR VGND sg13g2_decap_8
XFILLER_43_956 VPWR VGND sg13g2_decap_8
XFILLER_15_647 VPWR VGND sg13g2_decap_8
XFILLER_11_875 VPWR VGND sg13g2_decap_4
X_5921__315 VPWR VGND net315 sg13g2_tiehi
XFILLER_10_363 VPWR VGND sg13g2_fill_2
XFILLER_38_728 VPWR VGND sg13g2_decap_8
XFILLER_19_920 VPWR VGND sg13g2_decap_8
XFILLER_46_761 VPWR VGND sg13g2_decap_8
XFILLER_19_997 VPWR VGND sg13g2_decap_8
XFILLER_33_422 VPWR VGND sg13g2_fill_2
XFILLER_33_455 VPWR VGND sg13g2_fill_2
X_4840_ _1696_ VPWR _1718_ VGND _1685_ _1697_ sg13g2_o21ai_1
XFILLER_34_956 VPWR VGND sg13g2_decap_8
XFILLER_14_691 VPWR VGND sg13g2_decap_8
X_4771_ VGND VPWR _2542_ net451 _0234_ _1654_ sg13g2_a21oi_1
X_3722_ _0718_ VPWR _0731_ VGND _0711_ _0719_ sg13g2_o21ai_1
X_3653_ mydesign.pe_inputs\[61\] _0643_ _0663_ _0665_ _0666_ VPWR VGND sg13g2_and4_1
X_3584_ _0609_ _0599_ _0607_ VPWR VGND sg13g2_xnor2_1
X_5323_ net481 VPWR _2141_ VGND net758 _2140_ sg13g2_o21ai_1
X_5254_ _2082_ _2080_ _2084_ VPWR VGND sg13g2_xor2_1
X_4205_ _1147_ _1160_ _1161_ VPWR VGND sg13g2_nor2_1
X_5185_ _2019_ VPWR _2020_ VGND _2017_ _2018_ sg13g2_o21ai_1
X_5972__213 VPWR VGND net213 sg13g2_tiehi
X_4136_ VGND VPWR net561 _1094_ _0158_ _1095_ sg13g2_a21oi_1
XFILLER_3_1020 VPWR VGND sg13g2_decap_8
X_4067_ _1025_ VPWR _1038_ VGND _1024_ _1028_ sg13g2_o21ai_1
XFILLER_25_945 VPWR VGND sg13g2_decap_8
XFILLER_11_105 VPWR VGND sg13g2_decap_4
XFILLER_40_959 VPWR VGND sg13g2_decap_8
X_4969_ _1822_ _1815_ _1824_ VPWR VGND sg13g2_xor2_1
XFILLER_47_525 VPWR VGND sg13g2_decap_4
XFILLER_15_400 VPWR VGND sg13g2_fill_1
XFILLER_27_260 VPWR VGND sg13g2_fill_1
XFILLER_43_753 VPWR VGND sg13g2_decap_8
XFILLER_16_956 VPWR VGND sg13g2_decap_8
XFILLER_27_282 VPWR VGND sg13g2_decap_4
X_5949__259 VPWR VGND net259 sg13g2_tiehi
XFILLER_31_915 VPWR VGND sg13g2_decap_8
XFILLER_15_499 VPWR VGND sg13g2_fill_2
XFILLER_8_47 VPWR VGND sg13g2_fill_1
XFILLER_7_676 VPWR VGND sg13g2_decap_4
XFILLER_6_131 VPWR VGND sg13g2_decap_4
XFILLER_10_193 VPWR VGND sg13g2_fill_2
XFILLER_26_4 VPWR VGND sg13g2_decap_4
XFILLER_38_558 VPWR VGND sg13g2_fill_2
XFILLER_19_750 VPWR VGND sg13g2_fill_2
XFILLER_25_208 VPWR VGND sg13g2_fill_1
X_5941_ net275 VGND VPWR net957 mydesign.pe_inputs\[43\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_5872_ net29 VGND VPWR net1028 mydesign.pe_inputs\[58\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_4823_ _1700_ _1683_ _1702_ VPWR VGND sg13g2_xor2_1
XFILLER_21_458 VPWR VGND sg13g2_fill_2
X_4754_ _1645_ _1636_ _1644_ VPWR VGND sg13g2_xnor2_1
X_3705_ _0715_ mydesign.accum\[116\] _0714_ VPWR VGND sg13g2_xnor2_1
X_4685_ _1580_ mydesign.accum\[59\] _1577_ VPWR VGND sg13g2_xnor2_1
X_3636_ VPWR VGND mydesign.weights\[1\]\[22\] _0651_ net461 mydesign.weights\[1\]\[18\]
+ _0652_ net495 sg13g2_a221oi_1
X_3567_ _0591_ _0590_ _0593_ VPWR VGND sg13g2_xor2_1
XFILLER_1_808 VPWR VGND sg13g2_decap_8
X_5306_ _2132_ net695 _2131_ VPWR VGND sg13g2_nand2_1
X_5237_ _2066_ _2065_ _2054_ _2068_ VPWR VGND sg13g2_a21o_1
X_3498_ _0528_ net558 net455 _0517_ VPWR VGND sg13g2_and3_1
XFILLER_29_514 VPWR VGND sg13g2_fill_1
X_5168_ VGND VPWR _2527_ net494 _0280_ _2005_ sg13g2_a21oi_1
X_4119_ VGND VPWR net561 _1078_ _0157_ _1079_ sg13g2_a21oi_1
X_5099_ VGND VPWR net585 _1940_ _0275_ _1941_ sg13g2_a21oi_1
XFILLER_17_12 VPWR VGND sg13g2_fill_2
XFILLER_25_775 VPWR VGND sg13g2_decap_4
XFILLER_9_908 VPWR VGND sg13g2_decap_4
XFILLER_13_959 VPWR VGND sg13g2_decap_8
XFILLER_33_33 VPWR VGND sg13g2_fill_1
XFILLER_21_981 VPWR VGND sg13g2_decap_8
X_5801__149 VPWR VGND net149 sg13g2_tiehi
XFILLER_4_679 VPWR VGND sg13g2_fill_2
X_6116__108 VPWR VGND net108 sg13g2_tiehi
XFILLER_0_852 VPWR VGND sg13g2_decap_8
Xhold7 mydesign.inputs\[2\]\[5\] VPWR VGND net413 sg13g2_dlygate4sd3_1
XFILLER_48_867 VPWR VGND sg13g2_decap_8
XFILLER_43_572 VPWR VGND sg13g2_decap_4
XFILLER_12_970 VPWR VGND sg13g2_decap_8
Xhold418 mydesign.pe_inputs\[22\] VPWR VGND net1037 sg13g2_dlygate4sd3_1
XFILLER_7_462 VPWR VGND sg13g2_fill_2
Xhold407 _0259_ VPWR VGND net1026 sg13g2_dlygate4sd3_1
X_4470_ _1392_ _1393_ _0194_ VPWR VGND sg13g2_nor2_1
X_3421_ _0466_ _0464_ _0412_ _0463_ _0405_ VPWR VGND sg13g2_a22oi_1
Xhold429 mydesign.accum\[12\] VPWR VGND net1048 sg13g2_dlygate4sd3_1
XFILLER_48_1021 VPWR VGND sg13g2_decap_8
X_6140_ net264 VGND VPWR net932 mydesign.weights\[3\]\[14\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3352_ _2584_ _0402_ _0067_ VPWR VGND sg13g2_nor2_1
X_3283_ _2668_ net782 _2685_ _0038_ VPWR VGND sg13g2_mux2_1
X_6071_ net180 VGND VPWR _0297_ mydesign.pe_inputs\[9\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_5022_ _1874_ _1872_ _1873_ VPWR VGND sg13g2_nand2_1
XFILLER_38_311 VPWR VGND sg13g2_fill_1
XFILLER_38_355 VPWR VGND sg13g2_decap_4
XFILLER_17_0 VPWR VGND sg13g2_decap_8
XFILLER_26_506 VPWR VGND sg13g2_decap_8
X_5924_ net309 VGND VPWR _0150_ mydesign.pe_inputs\[46\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_5855_ net63 VGND VPWR _0081_ mydesign.pe_inputs\[61\] clknet_leaf_13_clk sg13g2_dfrbpq_2
XFILLER_21_222 VPWR VGND sg13g2_fill_1
XFILLER_21_233 VPWR VGND sg13g2_decap_4
XFILLER_22_756 VPWR VGND sg13g2_decap_4
X_4806_ _1685_ mydesign.pe_weights\[40\] mydesign.pe_inputs\[31\] VPWR VGND sg13g2_nand2_1
X_5786_ net165 VGND VPWR net663 mydesign.weights\[2\]\[19\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_4737_ VGND VPWR net567 _1628_ _0225_ _1629_ sg13g2_a21oi_1
X_4668_ _1564_ _1563_ _1555_ VPWR VGND sg13g2_nand2b_1
X_3619_ net630 VPWR _0638_ VGND net1059 net487 sg13g2_o21ai_1
X_4599_ VGND VPWR _1505_ _1506_ _1507_ net501 sg13g2_a21oi_1
X_5865__43 VPWR VGND net43 sg13g2_tiehi
XFILLER_29_322 VPWR VGND sg13g2_decap_8
XFILLER_44_43 VPWR VGND sg13g2_fill_2
XFILLER_25_550 VPWR VGND sg13g2_decap_8
XFILLER_44_65 VPWR VGND sg13g2_decap_4
XFILLER_13_745 VPWR VGND sg13g2_decap_4
XFILLER_12_299 VPWR VGND sg13g2_fill_1
XFILLER_48_664 VPWR VGND sg13g2_decap_8
X_3970_ _0947_ _0945_ _0946_ VPWR VGND sg13g2_nand2_1
X_5640_ _2429_ mydesign.pe_inputs\[6\] mydesign.pe_weights\[19\] VPWR VGND sg13g2_nand2_1
X_5571_ _2364_ mydesign.accum\[1\] mydesign.pe_inputs\[5\] net523 VPWR VGND sg13g2_and3_1
X_4522_ _1434_ _1416_ _1433_ VPWR VGND sg13g2_nand2_1
Xhold226 _1770_ VPWR VGND net845 sg13g2_dlygate4sd3_1
Xhold204 mydesign.weights\[3\]\[13\] VPWR VGND net823 sg13g2_dlygate4sd3_1
Xhold215 mydesign.out\[1\] VPWR VGND net834 sg13g2_dlygate4sd3_1
X_4453_ _1378_ _1358_ _1361_ _1377_ VPWR VGND sg13g2_and3_1
Xhold237 mydesign.pe_weights\[41\] VPWR VGND net856 sg13g2_dlygate4sd3_1
Xhold248 mydesign.compute_en VPWR VGND net867 sg13g2_dlygate4sd3_1
X_3404_ VGND VPWR _0441_ _0449_ _0071_ _0450_ sg13g2_a21oi_1
Xhold259 _0106_ VPWR VGND net878 sg13g2_dlygate4sd3_1
X_4384_ _1312_ _1310_ _1311_ VPWR VGND sg13g2_nand2_1
X_3335_ net544 net555 _0390_ VPWR VGND sg13g2_nor2b_2
X_6123_ net48 VGND VPWR _0349_ mydesign.weights\[1\]\[13\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_3266_ net616 VPWR _2676_ VGND net810 _2673_ sg13g2_o21ai_1
X_6054_ net242 VGND VPWR _0280_ mydesign.pe_inputs\[12\] clknet_leaf_29_clk sg13g2_dfrbpq_2
XFILLER_39_642 VPWR VGND sg13g2_decap_8
XFILLER_22_1024 VPWR VGND sg13g2_decap_4
X_5005_ _1857_ _1854_ _1858_ VPWR VGND sg13g2_xor2_1
XFILLER_39_664 VPWR VGND sg13g2_decap_4
X_3197_ net738 _2623_ net620 _2630_ VPWR VGND sg13g2_nand3_1
XFILLER_38_163 VPWR VGND sg13g2_fill_1
XFILLER_41_306 VPWR VGND sg13g2_decap_8
X_5907_ net340 VGND VPWR _0133_ mydesign.inputs\[0\]\[21\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5838_ net93 VGND VPWR _0064_ mydesign.cp\[2\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_5769_ _2513_ VPWR _0373_ VGND net602 _2511_ sg13g2_o21ai_1
X_5980__197 VPWR VGND net197 sg13g2_tiehi
XFILLER_30_56 VPWR VGND sg13g2_fill_2
XFILLER_2_914 VPWR VGND sg13g2_decap_8
XFILLER_2_903 VPWR VGND sg13g2_decap_8
XFILLER_49_439 VPWR VGND sg13g2_decap_4
X_6052__250 VPWR VGND net250 sg13g2_tiehi
XFILLER_29_196 VPWR VGND sg13g2_decap_8
XFILLER_45_667 VPWR VGND sg13g2_decap_8
XFILLER_44_188 VPWR VGND sg13g2_fill_1
XFILLER_41_895 VPWR VGND sg13g2_decap_8
XFILLER_9_557 VPWR VGND sg13g2_decap_4
XFILLER_45_1024 VPWR VGND sg13g2_decap_4
X_3120_ VPWR _2561_ net981 VGND sg13g2_inv_1
XFILLER_49_951 VPWR VGND sg13g2_decap_8
X_6031__334 VPWR VGND net334 sg13g2_tiehi
XFILLER_23_306 VPWR VGND sg13g2_decap_8
XFILLER_23_317 VPWR VGND sg13g2_fill_2
X_3953_ _0932_ net541 mydesign.weights\[3\]\[3\] net496 VPWR VGND sg13g2_and3_1
X_3884_ _0874_ _0855_ _0873_ VPWR VGND sg13g2_xnor2_1
X_5623_ _2413_ _2411_ _2412_ VPWR VGND sg13g2_nand2_1
X_5554_ net481 VPWR _2353_ VGND net592 net1055 sg13g2_o21ai_1
X_4505_ _1416_ _1417_ _1418_ VPWR VGND sg13g2_nor2b_1
X_5485_ _2288_ _2265_ _2287_ VPWR VGND sg13g2_nand2_1
X_4436_ VGND VPWR _1360_ _1361_ _1362_ net501 sg13g2_a21oi_1
Xfanout503 _2516_ net503 VPWR VGND sg13g2_buf_8
X_4367_ net473 VPWR _1297_ VGND net684 _1296_ sg13g2_o21ai_1
Xfanout514 net517 net514 VPWR VGND sg13g2_buf_8
Xfanout536 net1100 net536 VPWR VGND sg13g2_buf_8
Xfanout547 net548 net547 VPWR VGND sg13g2_buf_8
X_3318_ net1044 VPWR _0378_ VGND _2603_ net431 sg13g2_o21ai_1
Xfanout525 mydesign.pe_weights\[22\] net525 VPWR VGND sg13g2_buf_8
X_6106_ net228 VGND VPWR _0332_ mydesign.weights\[1\]\[16\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_4298_ _1239_ VPWR _1240_ VGND _1218_ _1220_ sg13g2_o21ai_1
Xfanout558 net562 net558 VPWR VGND sg13g2_buf_8
Xfanout569 net571 net569 VPWR VGND sg13g2_buf_8
X_6037_ net310 VGND VPWR _0263_ mydesign.accum\[43\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3249_ net2 _2666_ _2668_ VPWR VGND sg13g2_and2_1
XFILLER_42_637 VPWR VGND sg13g2_decap_4
XFILLER_26_188 VPWR VGND sg13g2_fill_2
XFILLER_10_501 VPWR VGND sg13g2_decap_8
XFILLER_10_512 VPWR VGND sg13g2_fill_1
XFILLER_22_383 VPWR VGND sg13g2_fill_2
XFILLER_46_943 VPWR VGND sg13g2_decap_8
XFILLER_17_100 VPWR VGND sg13g2_decap_8
XFILLER_17_155 VPWR VGND sg13g2_fill_2
XFILLER_14_851 VPWR VGND sg13g2_fill_2
XFILLER_41_692 VPWR VGND sg13g2_fill_1
XFILLER_40_180 VPWR VGND sg13g2_fill_2
XFILLER_12_1012 VPWR VGND sg13g2_decap_8
X_5959__239 VPWR VGND net239 sg13g2_tiehi
X_5270_ _2099_ _2097_ _2098_ VPWR VGND sg13g2_nand2_1
X_6139__280 VPWR VGND net280 sg13g2_tiehi
X_4221_ VGND VPWR _2571_ net447 _0164_ _1174_ sg13g2_a21oi_1
X_4152_ _1109_ _1108_ _1084_ _1111_ VPWR VGND sg13g2_a21o_1
X_4083_ net626 VPWR _1052_ VGND net489 _1051_ sg13g2_o21ai_1
XFILLER_37_910 VPWR VGND sg13g2_decap_8
X_3103_ VPWR _2544_ net1013 VGND sg13g2_inv_1
XFILLER_36_420 VPWR VGND sg13g2_fill_1
XFILLER_37_987 VPWR VGND sg13g2_decap_8
X_4985_ _1838_ _1835_ _1839_ VPWR VGND sg13g2_xor2_1
XFILLER_23_114 VPWR VGND sg13g2_decap_4
XFILLER_24_648 VPWR VGND sg13g2_fill_1
X_3936_ net459 VPWR _0917_ VGND mydesign.weights\[3\]\[9\] net547 sg13g2_o21ai_1
X_6107__224 VPWR VGND net224 sg13g2_tiehi
X_3867_ _0857_ mydesign.pe_inputs\[59\] _0789_ VPWR VGND sg13g2_nand2_1
X_5606_ _2397_ _2390_ _2396_ VPWR VGND sg13g2_nand2_1
X_3798_ mydesign.weights\[2\]\[18\] mydesign.weights\[2\]\[14\] net551 _0794_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_3_519 VPWR VGND sg13g2_decap_8
XFILLER_3_508 VPWR VGND sg13g2_fill_2
X_5537_ VPWR _2337_ _2336_ VGND sg13g2_inv_1
X_5468_ _2272_ _2253_ _2270_ VPWR VGND sg13g2_xnor2_1
X_5399_ VGND VPWR _2212_ _2211_ _2208_ sg13g2_or2_1
X_4419_ _1328_ VPWR _1345_ VGND _1327_ _1330_ sg13g2_o21ai_1
XFILLER_27_420 VPWR VGND sg13g2_fill_1
XFILLER_43_935 VPWR VGND sg13g2_decap_8
XFILLER_28_998 VPWR VGND sg13g2_decap_8
XFILLER_10_342 VPWR VGND sg13g2_fill_1
XFILLER_7_869 VPWR VGND sg13g2_decap_8
XFILLER_35_9 VPWR VGND sg13g2_fill_1
XFILLER_46_740 VPWR VGND sg13g2_decap_8
XFILLER_19_976 VPWR VGND sg13g2_decap_8
XFILLER_34_935 VPWR VGND sg13g2_decap_8
XFILLER_33_467 VPWR VGND sg13g2_fill_2
XFILLER_33_489 VPWR VGND sg13g2_fill_1
X_4770_ net637 VPWR _1654_ VGND mydesign.pe_weights\[26\] net452 sg13g2_o21ai_1
X_3721_ _0723_ _0727_ _0730_ VPWR VGND sg13g2_nor2_1
X_3652_ _0648_ net540 mydesign.accum\[113\] _0665_ VPWR VGND sg13g2_a21o_1
X_3583_ _0608_ _0599_ _0607_ VPWR VGND sg13g2_nand2_1
X_5322_ _2140_ net591 net522 mydesign.pe_weights\[24\] VPWR VGND sg13g2_and3_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_5253_ _2080_ _2082_ _2083_ VPWR VGND sg13g2_nor2_1
X_4204_ _1158_ _1156_ _1160_ VPWR VGND sg13g2_xor2_1
X_5184_ _2019_ _0395_ mydesign.inputs\[3\]\[15\] _2596_ mydesign.inputs\[3\]\[3\]
+ VPWR VGND sg13g2_a22oi_1
X_4135_ net468 VPWR _1095_ VGND net560 net964 sg13g2_o21ai_1
X_4066_ VGND VPWR _1023_ _1034_ _1037_ _1033_ sg13g2_a21oi_1
XFILLER_19_1018 VPWR VGND sg13g2_decap_8
XFILLER_40_938 VPWR VGND sg13g2_decap_8
X_4968_ _1815_ _1822_ _1823_ VPWR VGND sg13g2_nor2_1
X_4899_ _1769_ net1 _1768_ VPWR VGND sg13g2_nand2_2
XFILLER_20_640 VPWR VGND sg13g2_fill_1
X_3919_ _0906_ net835 _0905_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_684 VPWR VGND sg13g2_fill_1
XFILLER_4_828 VPWR VGND sg13g2_decap_4
XFILLER_16_935 VPWR VGND sg13g2_decap_8
XFILLER_43_732 VPWR VGND sg13g2_decap_8
XFILLER_11_640 VPWR VGND sg13g2_fill_2
XFILLER_10_161 VPWR VGND sg13g2_decap_8
XFILLER_6_143 VPWR VGND sg13g2_decap_8
XFILLER_3_861 VPWR VGND sg13g2_fill_2
XFILLER_19_740 VPWR VGND sg13g2_fill_2
XFILLER_19_784 VPWR VGND sg13g2_fill_2
X_5940_ net277 VGND VPWR _0166_ mydesign.pe_inputs\[42\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_5871_ net31 VGND VPWR net1016 mydesign.pe_inputs\[57\] clknet_leaf_42_clk sg13g2_dfrbpq_2
XFILLER_22_905 VPWR VGND sg13g2_decap_4
XFILLER_33_242 VPWR VGND sg13g2_fill_2
XFILLER_21_415 VPWR VGND sg13g2_fill_2
X_4822_ _1700_ _1683_ _1701_ VPWR VGND sg13g2_nor2b_1
X_4753_ _1643_ net941 _1644_ VPWR VGND sg13g2_xor2_1
X_3704_ mydesign.pe_inputs\[61\] _0658_ _0714_ VPWR VGND sg13g2_and2_1
X_4684_ mydesign.accum\[59\] _1577_ _1579_ VPWR VGND sg13g2_nor2b_1
X_3635_ _0651_ net545 net556 mydesign.weights\[1\]\[14\] VPWR VGND sg13g2_and3_1
X_3566_ _0592_ _0591_ _0590_ VPWR VGND sg13g2_nand2b_1
X_3497_ VGND VPWR _2575_ net485 _0087_ _0527_ sg13g2_a21oi_1
X_5305_ VGND VPWR net611 _2640_ _2131_ net608 sg13g2_a21oi_1
X_5236_ _2065_ _2066_ _2054_ _2067_ VPWR VGND sg13g2_nand3_1
XFILLER_25_1022 VPWR VGND sg13g2_decap_8
X_5167_ net625 VPWR _2005_ VGND net489 _2004_ sg13g2_o21ai_1
XFILLER_29_537 VPWR VGND sg13g2_decap_8
X_4118_ net468 VPWR _1079_ VGND net561 net896 sg13g2_o21ai_1
X_5098_ net475 VPWR _1941_ VGND net585 net864 sg13g2_o21ai_1
X_4049_ VGND VPWR net565 _1020_ _0145_ _1021_ sg13g2_a21oi_1
XFILLER_37_592 VPWR VGND sg13g2_decap_8
XFILLER_37_581 VPWR VGND sg13g2_decap_4
XFILLER_17_68 VPWR VGND sg13g2_decap_8
XFILLER_13_938 VPWR VGND sg13g2_decap_8
XFILLER_33_23 VPWR VGND sg13g2_fill_1
XFILLER_12_459 VPWR VGND sg13g2_decap_8
XFILLER_21_960 VPWR VGND sg13g2_decap_8
XFILLER_0_831 VPWR VGND sg13g2_decap_8
XFILLER_48_846 VPWR VGND sg13g2_decap_8
Xhold8 mydesign.inputs\[2\]\[12\] VPWR VGND net414 sg13g2_dlygate4sd3_1
X_5990__166 VPWR VGND net166 sg13g2_tiehi
XFILLER_28_581 VPWR VGND sg13g2_fill_2
XFILLER_43_562 VPWR VGND sg13g2_fill_1
XFILLER_16_776 VPWR VGND sg13g2_decap_8
XFILLER_31_702 VPWR VGND sg13g2_decap_4
Xhold408 mydesign.pe_inputs\[58\] VPWR VGND net1027 sg13g2_dlygate4sd3_1
XFILLER_48_1000 VPWR VGND sg13g2_decap_8
X_3420_ net513 mydesign.accum\[101\] mydesign.accum\[69\] mydesign.accum\[37\] mydesign.accum\[5\]
+ net506 _0465_ VPWR VGND sg13g2_mux4_1
Xhold419 mydesign.accum\[10\] VPWR VGND net1038 sg13g2_dlygate4sd3_1
X_3351_ VGND VPWR _2585_ _0400_ _0066_ _0402_ sg13g2_a21oi_1
X_6070_ net186 VGND VPWR net1099 mydesign.pe_inputs\[8\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_3282_ _2667_ net796 _2685_ _0037_ VPWR VGND sg13g2_mux2_1
XFILLER_39_824 VPWR VGND sg13g2_fill_2
X_5021_ mydesign.pe_inputs\[27\] mydesign.pe_weights\[39\] mydesign.accum\[46\] _1873_
+ VPWR VGND sg13g2_a21o_1
XFILLER_39_879 VPWR VGND sg13g2_decap_8
XFILLER_38_378 VPWR VGND sg13g2_fill_1
XFILLER_0_1013 VPWR VGND sg13g2_decap_8
X_5923_ net311 VGND VPWR _0149_ mydesign.pe_inputs\[45\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_5854_ net65 VGND VPWR _0080_ mydesign.pe_inputs\[60\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_4805_ _1675_ VPWR _1684_ VGND _1668_ _1676_ sg13g2_o21ai_1
X_5785_ net167 VGND VPWR _0011_ mydesign.weights\[2\]\[18\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_4736_ net469 VPWR _1629_ VGND net567 net840 sg13g2_o21ai_1
X_4667_ _1563_ _1545_ _1561_ VPWR VGND sg13g2_xnor2_1
X_3618_ VGND VPWR _2581_ net490 _0098_ _0637_ sg13g2_a21oi_1
X_4598_ _1504_ VPWR _1506_ VGND _1491_ _1494_ sg13g2_o21ai_1
X_3549_ VGND VPWR _0574_ _0575_ _0576_ net499 sg13g2_a21oi_1
XFILLER_0_116 VPWR VGND sg13g2_fill_2
X_5800__150 VPWR VGND net150 sg13g2_tiehi
XFILLER_0_149 VPWR VGND sg13g2_decap_4
X_5219_ VGND VPWR net563 _2049_ _0286_ _2050_ sg13g2_a21oi_1
XFILLER_45_849 VPWR VGND sg13g2_decap_8
XFILLER_44_55 VPWR VGND sg13g2_fill_1
XFILLER_21_790 VPWR VGND sg13g2_decap_4
XFILLER_5_901 VPWR VGND sg13g2_decap_8
XFILLER_4_444 VPWR VGND sg13g2_fill_2
XFILLER_0_650 VPWR VGND sg13g2_decap_8
XFILLER_48_643 VPWR VGND sg13g2_decap_8
XFILLER_0_694 VPWR VGND sg13g2_decap_4
XFILLER_36_849 VPWR VGND sg13g2_fill_1
XFILLER_43_370 VPWR VGND sg13g2_decap_8
XFILLER_15_1021 VPWR VGND sg13g2_decap_8
X_5570_ _2363_ mydesign.pe_inputs\[4\] mydesign.pe_weights\[17\] VPWR VGND sg13g2_nand2_1
X_4521_ _1433_ _1423_ _1432_ VPWR VGND sg13g2_xnor2_1
X_5997__106 VPWR VGND net106 sg13g2_tiehi
Xhold205 _2507_ VPWR VGND net824 sg13g2_dlygate4sd3_1
X_4452_ _1375_ _1354_ _1377_ VPWR VGND sg13g2_xor2_1
Xhold216 mydesign.accum\[111\] VPWR VGND net835 sg13g2_dlygate4sd3_1
Xhold227 _0248_ VPWR VGND net846 sg13g2_dlygate4sd3_1
Xhold249 mydesign.accum\[75\] VPWR VGND net868 sg13g2_dlygate4sd3_1
X_3403_ net627 VPWR _0450_ VGND net1078 net430 sg13g2_o21ai_1
Xhold238 _0233_ VPWR VGND net857 sg13g2_dlygate4sd3_1
X_4383_ net534 mydesign.pe_weights\[54\] mydesign.accum\[74\] _1311_ VPWR VGND sg13g2_a21o_1
X_3334_ _0062_ net613 _0388_ _0389_ VPWR VGND sg13g2_and3_1
X_6122_ net56 VGND VPWR _0348_ mydesign.weights\[1\]\[12\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_6053_ net246 VGND VPWR _0279_ mydesign.accum\[39\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_3265_ VGND VPWR _2519_ _2673_ _0030_ _2675_ sg13g2_a21oi_1
X_5938__281 VPWR VGND net281 sg13g2_tiehi
XFILLER_22_1003 VPWR VGND sg13g2_decap_8
X_5004_ _1857_ _1855_ _1856_ VPWR VGND sg13g2_nand2_1
X_3196_ _2628_ VPWR _0007_ VGND _2623_ net600 sg13g2_o21ai_1
XFILLER_38_131 VPWR VGND sg13g2_fill_1
X_5969__219 VPWR VGND net219 sg13g2_tiehi
X_5906_ net341 VGND VPWR _0132_ mydesign.inputs\[0\]\[20\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5837_ net95 VGND VPWR _0063_ mydesign.cp\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_10_727 VPWR VGND sg13g2_fill_2
XFILLER_10_749 VPWR VGND sg13g2_fill_1
X_5768_ _2513_ net693 _2511_ VPWR VGND sg13g2_nand2_1
X_4719_ VGND VPWR net567 _1611_ _0224_ _1612_ sg13g2_a21oi_1
X_5699_ net725 _2476_ net613 _2477_ VPWR VGND sg13g2_nand3_1
XFILLER_1_425 VPWR VGND sg13g2_decap_4
XFILLER_17_304 VPWR VGND sg13g2_fill_1
XFILLER_45_646 VPWR VGND sg13g2_decap_8
XFILLER_44_112 VPWR VGND sg13g2_fill_2
XFILLER_38_1021 VPWR VGND sg13g2_decap_8
XFILLER_25_370 VPWR VGND sg13g2_fill_1
XFILLER_32_318 VPWR VGND sg13g2_fill_2
XFILLER_41_874 VPWR VGND sg13g2_decap_8
XFILLER_5_753 VPWR VGND sg13g2_decap_4
XFILLER_45_1003 VPWR VGND sg13g2_decap_8
XFILLER_49_930 VPWR VGND sg13g2_decap_8
XFILLER_1_992 VPWR VGND sg13g2_decap_8
XFILLER_36_635 VPWR VGND sg13g2_fill_2
XFILLER_36_668 VPWR VGND sg13g2_fill_2
XFILLER_17_882 VPWR VGND sg13g2_fill_1
XFILLER_17_893 VPWR VGND sg13g2_fill_1
X_3952_ _0931_ mydesign.weights\[3\]\[15\] _2586_ _0394_ VPWR VGND sg13g2_and3_1
X_3883_ _0873_ _0872_ _0871_ VPWR VGND sg13g2_nand2b_1
X_5622_ mydesign.pe_weights\[17\] net519 mydesign.accum\[4\] _2412_ VPWR VGND sg13g2_a21o_1
X_5553_ _2351_ _2348_ _2352_ VPWR VGND sg13g2_xor2_1
X_4504_ _1415_ VPWR _1417_ VGND _1413_ _1414_ sg13g2_o21ai_1
X_5484_ _2285_ _2278_ _2287_ VPWR VGND sg13g2_xor2_1
X_4435_ _1359_ VPWR _1361_ VGND _1339_ _1341_ sg13g2_o21ai_1
X_4366_ net501 _2559_ _2563_ _1296_ VPWR VGND sg13g2_nor3_1
Xfanout504 net510 net504 VPWR VGND sg13g2_buf_8
Xfanout515 net516 net515 VPWR VGND sg13g2_buf_8
Xfanout548 net553 net548 VPWR VGND sg13g2_buf_1
X_3317_ VGND VPWR net842 _0376_ _0057_ _0377_ sg13g2_a21oi_1
Xfanout537 net1067 net537 VPWR VGND sg13g2_buf_8
X_6105_ net236 VGND VPWR net410 mydesign.accum\[7\] clknet_leaf_39_clk sg13g2_dfrbpq_1
Xfanout526 net1097 net526 VPWR VGND sg13g2_buf_8
X_4297_ _1238_ _1230_ _1239_ VPWR VGND sg13g2_xor2_1
Xfanout559 net562 net559 VPWR VGND sg13g2_buf_1
XFILLER_39_451 VPWR VGND sg13g2_fill_2
X_6036_ net314 VGND VPWR net922 mydesign.accum\[42\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3248_ net794 _2667_ _2659_ _0021_ VPWR VGND sg13g2_mux2_1
XFILLER_39_473 VPWR VGND sg13g2_fill_1
X_3179_ _2616_ net752 net623 VPWR VGND sg13g2_nand2_1
XFILLER_23_841 VPWR VGND sg13g2_fill_1
XFILLER_41_12 VPWR VGND sg13g2_decap_8
XFILLER_1_222 VPWR VGND sg13g2_fill_2
XFILLER_2_789 VPWR VGND sg13g2_fill_2
XFILLER_1_288 VPWR VGND sg13g2_fill_1
XFILLER_2_28 VPWR VGND sg13g2_fill_2
XFILLER_46_922 VPWR VGND sg13g2_decap_8
XFILLER_18_646 VPWR VGND sg13g2_decap_8
XFILLER_46_999 VPWR VGND sg13g2_decap_8
XFILLER_45_487 VPWR VGND sg13g2_fill_2
XFILLER_14_830 VPWR VGND sg13g2_fill_1
XFILLER_14_841 VPWR VGND sg13g2_fill_1
XFILLER_32_137 VPWR VGND sg13g2_fill_2
XFILLER_41_682 VPWR VGND sg13g2_fill_1
XFILLER_40_170 VPWR VGND sg13g2_fill_2
XFILLER_5_583 VPWR VGND sg13g2_fill_2
XFILLER_5_561 VPWR VGND sg13g2_fill_1
X_4220_ net631 VPWR _1174_ VGND net1050 net447 sg13g2_o21ai_1
X_4151_ _1108_ _1109_ _1084_ _1110_ VPWR VGND sg13g2_nand3_1
X_4082_ _1048_ VPWR _1051_ VGND net542 _1050_ sg13g2_o21ai_1
X_6085__28 VPWR VGND net28 sg13g2_tiehi
X_3102_ VPWR _2543_ net856 VGND sg13g2_inv_1
XFILLER_37_966 VPWR VGND sg13g2_decap_8
X_4984_ _1838_ _1836_ _1837_ VPWR VGND sg13g2_nand2_1
X_3935_ net497 mydesign.weights\[3\]\[5\] _0916_ VPWR VGND sg13g2_nor2_1
XFILLER_20_833 VPWR VGND sg13g2_decap_8
XFILLER_32_682 VPWR VGND sg13g2_fill_1
X_5605_ _2396_ _2391_ _2395_ VPWR VGND sg13g2_xnor2_1
X_3866_ _0845_ VPWR _0856_ VGND _0820_ _0843_ sg13g2_o21ai_1
X_3797_ _0791_ _0792_ net459 _0793_ VPWR VGND sg13g2_nand3_1
XFILLER_20_888 VPWR VGND sg13g2_fill_2
X_5536_ _2318_ VPWR _2336_ VGND _2316_ _2319_ sg13g2_o21ai_1
X_5467_ _2271_ _2253_ _2270_ VPWR VGND sg13g2_nand2_1
X_4418_ _1344_ mydesign.pe_weights\[53\] mydesign.pe_inputs\[43\] VPWR VGND sg13g2_nand2_1
X_5398_ _2211_ _2209_ _2210_ VPWR VGND sg13g2_nand2_1
X_4349_ VGND VPWR net580 _1286_ _0179_ _1287_ sg13g2_a21oi_1
XFILLER_47_719 VPWR VGND sg13g2_decap_8
XFILLER_39_270 VPWR VGND sg13g2_decap_8
X_6019_ net390 VGND VPWR _0245_ mydesign.inputs\[3\]\[5\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_27_454 VPWR VGND sg13g2_decap_4
XFILLER_28_977 VPWR VGND sg13g2_decap_8
XFILLER_43_914 VPWR VGND sg13g2_decap_8
XFILLER_15_605 VPWR VGND sg13g2_fill_1
XFILLER_27_487 VPWR VGND sg13g2_decap_8
XFILLER_35_1013 VPWR VGND sg13g2_decap_8
XFILLER_2_564 VPWR VGND sg13g2_fill_2
XFILLER_42_1017 VPWR VGND sg13g2_decap_8
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_37_207 VPWR VGND sg13g2_decap_4
XFILLER_37_218 VPWR VGND sg13g2_decap_4
XFILLER_19_955 VPWR VGND sg13g2_decap_8
XFILLER_46_796 VPWR VGND sg13g2_decap_8
XFILLER_45_240 VPWR VGND sg13g2_decap_8
XFILLER_34_914 VPWR VGND sg13g2_decap_8
XFILLER_33_424 VPWR VGND sg13g2_fill_1
X_3720_ VGND VPWR net577 _0728_ _0108_ _0729_ sg13g2_a21oi_1
Xclkbuf_leaf_40_clk clknet_3_4__leaf_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
X_3651_ VPWR _0664_ _0663_ VGND sg13g2_inv_1
X_3582_ _0605_ _0604_ _0607_ VPWR VGND sg13g2_xor2_1
X_5321_ VGND VPWR _2525_ net449 _0299_ _2139_ sg13g2_a21oi_1
X_5252_ _2082_ mydesign.accum\[28\] _2081_ VPWR VGND sg13g2_xnor2_1
X_4203_ _1159_ _1156_ _1158_ VPWR VGND sg13g2_nand2b_1
X_5183_ net459 VPWR _2018_ VGND net549 mydesign.inputs\[3\]\[11\] sg13g2_o21ai_1
X_4134_ _1093_ _1076_ _1094_ VPWR VGND sg13g2_xor2_1
XFILLER_3_60 VPWR VGND sg13g2_fill_2
XFILLER_28_229 VPWR VGND sg13g2_fill_2
XFILLER_37_730 VPWR VGND sg13g2_fill_1
X_4065_ VGND VPWR net566 _1035_ _0146_ _1036_ sg13g2_a21oi_1
XFILLER_40_917 VPWR VGND sg13g2_decap_8
X_4967_ _1820_ _1799_ _1822_ VPWR VGND sg13g2_xor2_1
XFILLER_33_980 VPWR VGND sg13g2_decap_8
X_5827__115 VPWR VGND net115 sg13g2_tiehi
X_4898_ VGND VPWR _2605_ _1768_ _2688_ _2664_ sg13g2_a21oi_2
Xclkbuf_leaf_31_clk clknet_3_6__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
X_3918_ _0894_ VPWR _0905_ VGND _0893_ _0896_ sg13g2_o21ai_1
X_3849_ mydesign.pe_inputs\[56\] _0804_ mydesign.accum\[107\] _0840_ VPWR VGND sg13g2_nand3_1
XFILLER_22_58 VPWR VGND sg13g2_fill_1
X_5519_ _2317_ _2319_ _2320_ VPWR VGND sg13g2_nor2_1
XFILLER_3_328 VPWR VGND sg13g2_fill_2
XFILLER_47_55 VPWR VGND sg13g2_fill_2
XFILLER_43_711 VPWR VGND sg13g2_decap_8
XFILLER_43_788 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_22_clk clknet_3_6__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_6_100 VPWR VGND sg13g2_fill_2
XFILLER_2_361 VPWR VGND sg13g2_decap_8
XFILLER_33_7 VPWR VGND sg13g2_decap_8
X_5870_ net33 VGND VPWR net1074 mydesign.pe_inputs\[56\] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_4821_ _1700_ _1684_ _1698_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_928 VPWR VGND sg13g2_fill_1
XFILLER_34_799 VPWR VGND sg13g2_fill_1
XFILLER_21_449 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_13_clk clknet_3_2__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_4752_ _1632_ VPWR _1643_ VGND _1631_ _1634_ sg13g2_o21ai_1
X_3703_ _0713_ mydesign.pe_inputs\[62\] _0653_ VPWR VGND sg13g2_nand2_1
X_4683_ net535 _1521_ mydesign.accum\[59\] _1578_ VPWR VGND sg13g2_nand3_1
XFILLER_30_983 VPWR VGND sg13g2_decap_8
X_3634_ mydesign.weights\[1\]\[10\] net460 net498 _0650_ VPWR VGND sg13g2_nand3_1
X_5904__345 VPWR VGND net345 sg13g2_tiehi
X_3565_ _0568_ VPWR _0591_ VGND _0557_ _0569_ sg13g2_o21ai_1
X_3496_ net624 VPWR _0527_ VGND net484 _0526_ sg13g2_o21ai_1
X_5304_ _2130_ net611 _2640_ VPWR VGND sg13g2_nand2_2
X_5235_ _2064_ _2063_ _2040_ _2066_ VPWR VGND sg13g2_a21o_1
XFILLER_25_1001 VPWR VGND sg13g2_decap_8
X_5166_ _2001_ _2002_ _2003_ _2004_ VPWR VGND sg13g2_or3_1
X_4117_ VGND VPWR _1078_ _1077_ _1076_ sg13g2_or2_1
X_5097_ _1938_ _1921_ _1940_ VPWR VGND sg13g2_xor2_1
XFILLER_17_14 VPWR VGND sg13g2_fill_1
X_4048_ net464 VPWR _1021_ VGND net565 net968 sg13g2_o21ai_1
X_5999_ net98 VGND VPWR _0225_ mydesign.accum\[61\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_25_788 VPWR VGND sg13g2_fill_1
X_5948__261 VPWR VGND net261 sg13g2_tiehi
XFILLER_32_1027 VPWR VGND sg13g2_fill_2
XFILLER_4_637 VPWR VGND sg13g2_fill_1
XFILLER_0_810 VPWR VGND sg13g2_decap_8
XFILLER_48_825 VPWR VGND sg13g2_decap_8
XFILLER_0_887 VPWR VGND sg13g2_decap_8
Xhold9 _0076_ VPWR VGND net415 sg13g2_dlygate4sd3_1
XFILLER_47_368 VPWR VGND sg13g2_decap_4
XFILLER_28_593 VPWR VGND sg13g2_fill_2
XFILLER_30_202 VPWR VGND sg13g2_fill_2
XFILLER_30_257 VPWR VGND sg13g2_fill_1
XFILLER_11_471 VPWR VGND sg13g2_fill_2
XFILLER_8_987 VPWR VGND sg13g2_decap_8
Xhold409 _0098_ VPWR VGND net1028 sg13g2_dlygate4sd3_1
X_3350_ net618 VPWR _0402_ VGND _2585_ _0400_ sg13g2_o21ai_1
X_3281_ _2685_ _2655_ _2684_ VPWR VGND sg13g2_nand2_2
X_5020_ net531 mydesign.pe_inputs\[27\] mydesign.accum\[46\] _1872_ VPWR VGND sg13g2_nand3_1
XFILLER_39_814 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_2_clk clknet_3_1__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
X_6034__322 VPWR VGND net322 sg13g2_tiehi
X_5817__125 VPWR VGND net125 sg13g2_tiehi
XFILLER_38_335 VPWR VGND sg13g2_fill_1
XFILLER_47_880 VPWR VGND sg13g2_decap_8
X_5922_ net313 VGND VPWR _0148_ mydesign.pe_inputs\[44\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_5853_ net66 VGND VPWR net653 mydesign.inputs\[2\]\[15\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_5784_ net169 VGND VPWR net676 mydesign.weights\[2\]\[17\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_4804_ _1679_ VPWR _1683_ VGND _1665_ _1680_ sg13g2_o21ai_1
X_4735_ _1628_ _1613_ _1627_ VPWR VGND sg13g2_xnor2_1
X_5824__118 VPWR VGND net118 sg13g2_tiehi
X_4666_ _1562_ _1561_ _1545_ VPWR VGND sg13g2_nand2b_1
X_4597_ _1491_ _1494_ _1504_ _1505_ VPWR VGND sg13g2_or3_1
X_3617_ net630 VPWR _0637_ VGND mydesign.pe_inputs\[62\] net487 sg13g2_o21ai_1
X_3548_ _0553_ _0551_ _0573_ _0575_ VPWR VGND sg13g2_a21o_1
X_3479_ net609 _0513_ _0083_ VPWR VGND sg13g2_nor2_1
X_6115__132 VPWR VGND net132 sg13g2_tiehi
X_5218_ net466 VPWR _2050_ VGND net563 net923 sg13g2_o21ai_1
X_5149_ _1975_ _1978_ _1988_ _1989_ VPWR VGND sg13g2_nor3_1
XFILLER_45_828 VPWR VGND sg13g2_decap_8
XFILLER_44_349 VPWR VGND sg13g2_fill_2
XFILLER_5_979 VPWR VGND sg13g2_decap_8
XFILLER_48_622 VPWR VGND sg13g2_decap_8
X_5775__183 VPWR VGND net183 sg13g2_tiehi
XFILLER_48_699 VPWR VGND sg13g2_decap_8
XFILLER_18_90 VPWR VGND sg13g2_fill_1
XFILLER_44_883 VPWR VGND sg13g2_decap_8
XFILLER_15_1000 VPWR VGND sg13g2_decap_8
XFILLER_31_588 VPWR VGND sg13g2_decap_4
X_4520_ _1429_ _1413_ _1432_ VPWR VGND sg13g2_xor2_1
XFILLER_11_290 VPWR VGND sg13g2_fill_2
Xhold217 mydesign.pe_inputs\[45\] VPWR VGND net836 sg13g2_dlygate4sd3_1
Xhold206 _0365_ VPWR VGND net825 sg13g2_dlygate4sd3_1
X_4451_ _1354_ _1375_ _1376_ VPWR VGND sg13g2_nor2b_1
Xhold228 mydesign.accum\[98\] VPWR VGND net847 sg13g2_dlygate4sd3_1
Xhold239 mydesign.weights\[3\]\[9\] VPWR VGND net858 sg13g2_dlygate4sd3_1
X_3402_ VPWR VGND _0412_ _0448_ _0443_ net456 _0449_ _0442_ sg13g2_a221oi_1
XFILLER_4_990 VPWR VGND sg13g2_decap_8
X_4382_ mydesign.pe_weights\[54\] net534 mydesign.accum\[74\] _1310_ VPWR VGND sg13g2_nand3_1
X_6121_ net64 VGND VPWR _0347_ mydesign.weights\[1\]\[11\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3333_ _0387_ VPWR _0389_ VGND net548 net454 sg13g2_o21ai_1
X_6052_ net250 VGND VPWR _0278_ mydesign.accum\[38\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_3264_ net616 VPWR _2675_ VGND net807 _2673_ sg13g2_o21ai_1
X_5003_ mydesign.pe_inputs\[26\] net531 mydesign.accum\[45\] _1856_ VPWR VGND sg13g2_a21o_1
X_3195_ _2629_ net3 net620 VPWR VGND sg13g2_nand2_2
XFILLER_26_316 VPWR VGND sg13g2_fill_2
XFILLER_42_809 VPWR VGND sg13g2_fill_2
X_5905_ net343 VGND VPWR _0131_ mydesign.accum\[111\] clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_35_894 VPWR VGND sg13g2_decap_8
XFILLER_22_544 VPWR VGND sg13g2_decap_8
XFILLER_34_382 VPWR VGND sg13g2_fill_2
X_5836_ net97 VGND VPWR _0062_ mydesign.cp\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_2
X_5767_ _2512_ VPWR _0372_ VGND net604 _2511_ sg13g2_o21ai_1
X_5698_ net610 _2656_ mydesign.load_counter\[3\] _2476_ VPWR VGND sg13g2_nand3_1
X_4718_ net467 VPWR _1612_ VGND net567 net866 sg13g2_o21ai_1
X_4649_ _1521_ mydesign.pe_weights\[45\] mydesign.accum\[57\] _1546_ VPWR VGND sg13g2_a21o_1
XFILLER_2_938 VPWR VGND sg13g2_fill_2
XFILLER_49_419 VPWR VGND sg13g2_decap_4
XFILLER_49_408 VPWR VGND sg13g2_fill_2
XFILLER_7_1009 VPWR VGND sg13g2_decap_8
XFILLER_29_132 VPWR VGND sg13g2_fill_1
XFILLER_45_625 VPWR VGND sg13g2_decap_8
XFILLER_17_316 VPWR VGND sg13g2_fill_1
XFILLER_44_135 VPWR VGND sg13g2_decap_8
XFILLER_44_124 VPWR VGND sg13g2_fill_2
XFILLER_44_179 VPWR VGND sg13g2_decap_8
XFILLER_38_1000 VPWR VGND sg13g2_decap_8
XFILLER_41_853 VPWR VGND sg13g2_decap_8
XFILLER_9_515 VPWR VGND sg13g2_decap_8
XFILLER_5_765 VPWR VGND sg13g2_fill_1
XFILLER_1_971 VPWR VGND sg13g2_decap_8
XFILLER_49_986 VPWR VGND sg13g2_decap_8
XFILLER_48_485 VPWR VGND sg13g2_fill_1
X_5814__128 VPWR VGND net128 sg13g2_tiehi
X_3951_ VGND VPWR _0928_ _0929_ _0930_ _0397_ sg13g2_a21oi_1
XFILLER_35_157 VPWR VGND sg13g2_fill_1
XFILLER_44_680 VPWR VGND sg13g2_decap_8
XFILLER_16_371 VPWR VGND sg13g2_fill_1
XFILLER_32_831 VPWR VGND sg13g2_fill_1
X_3882_ _0872_ _0869_ _0870_ VPWR VGND sg13g2_nand2b_1
XFILLER_31_341 VPWR VGND sg13g2_decap_8
X_5621_ net519 mydesign.pe_weights\[17\] mydesign.accum\[4\] _2411_ VPWR VGND sg13g2_nand3_1
X_5552_ _2351_ _2339_ _2350_ VPWR VGND sg13g2_xnor2_1
X_4503_ _1413_ _1414_ _1415_ _1416_ VPWR VGND sg13g2_nor3_1
X_5483_ _2278_ _2285_ _2286_ VPWR VGND sg13g2_nor2_1
X_4434_ _1339_ _1341_ _1359_ _1360_ VPWR VGND sg13g2_or3_1
X_4365_ VGND VPWR _2533_ net493 _0187_ _1295_ sg13g2_a21oi_1
Xfanout505 net510 net505 VPWR VGND sg13g2_buf_8
Xfanout527 mydesign.pe_weights\[27\] net527 VPWR VGND sg13g2_buf_8
X_3316_ net613 VPWR _0377_ VGND net842 _2600_ sg13g2_o21ai_1
X_6104_ net244 VGND VPWR _0330_ mydesign.accum\[6\] clknet_leaf_37_clk sg13g2_dfrbpq_2
Xfanout538 net1092 net538 VPWR VGND sg13g2_buf_8
Xfanout516 net517 net516 VPWR VGND sg13g2_buf_8
X_4296_ _1238_ _1231_ _1236_ VPWR VGND sg13g2_xnor2_1
Xfanout549 net552 net549 VPWR VGND sg13g2_buf_8
X_6035_ net318 VGND VPWR net950 mydesign.accum\[41\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3247_ net1 _2666_ _2667_ VPWR VGND sg13g2_and2_1
X_3178_ _2615_ net4 net432 VPWR VGND sg13g2_nand2_1
XFILLER_27_658 VPWR VGND sg13g2_fill_2
XFILLER_22_385 VPWR VGND sg13g2_fill_1
X_5819_ net123 VGND VPWR _0045_ mydesign.inputs\[0\]\[12\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_10_547 VPWR VGND sg13g2_decap_8
XFILLER_46_901 VPWR VGND sg13g2_decap_8
XFILLER_46_978 VPWR VGND sg13g2_decap_8
XFILLER_32_105 VPWR VGND sg13g2_fill_1
XFILLER_32_116 VPWR VGND sg13g2_decap_4
XFILLER_13_341 VPWR VGND sg13g2_fill_2
XFILLER_14_853 VPWR VGND sg13g2_fill_1
XFILLER_13_374 VPWR VGND sg13g2_fill_2
XFILLER_40_182 VPWR VGND sg13g2_fill_1
X_4150_ _1100_ VPWR _1109_ VGND _1106_ _1107_ sg13g2_o21ai_1
X_3101_ VPWR _2542_ net813 VGND sg13g2_inv_1
X_4081_ VPWR VGND mydesign.inputs\[1\]\[21\] _1049_ net461 mydesign.inputs\[1\]\[17\]
+ _1050_ net495 sg13g2_a221oi_1
XFILLER_49_783 VPWR VGND sg13g2_decap_8
XFILLER_48_293 VPWR VGND sg13g2_decap_8
XFILLER_37_945 VPWR VGND sg13g2_decap_8
X_4983_ mydesign.pe_inputs\[25\] net531 mydesign.accum\[44\] _1837_ VPWR VGND sg13g2_a21o_1
X_3934_ VGND VPWR net433 _0914_ _0136_ _0915_ sg13g2_a21oi_1
X_3865_ _0851_ VPWR _0855_ VGND _0834_ _0852_ sg13g2_o21ai_1
X_5604_ _2392_ _2394_ _2395_ VPWR VGND sg13g2_nor2_1
XFILLER_31_182 VPWR VGND sg13g2_decap_4
X_3796_ VGND VPWR _0792_ mydesign.weights\[2\]\[10\] net549 sg13g2_or2_1
XFILLER_20_878 VPWR VGND sg13g2_fill_2
X_5535_ _2335_ _2334_ _2333_ VPWR VGND sg13g2_nand2b_1
X_5466_ _2270_ _2260_ _2269_ VPWR VGND sg13g2_xnor2_1
X_4417_ VGND VPWR net576 _1342_ _0191_ _1343_ sg13g2_a21oi_1
X_5397_ net527 mydesign.pe_inputs\[14\] mydesign.accum\[21\] _2210_ VPWR VGND sg13g2_a21o_1
X_4348_ net479 VPWR _1287_ VGND net579 net865 sg13g2_o21ai_1
X_4279_ _1222_ _1199_ _1221_ VPWR VGND sg13g2_nand2_1
X_6018_ net394 VGND VPWR _0244_ mydesign.inputs\[3\]\[4\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_27_411 VPWR VGND sg13g2_decap_8
XFILLER_28_956 VPWR VGND sg13g2_decap_8
XFILLER_10_333 VPWR VGND sg13g2_decap_8
XFILLER_6_359 VPWR VGND sg13g2_fill_2
XFILLER_10_399 VPWR VGND sg13g2_fill_2
X_5958__241 VPWR VGND net241 sg13g2_tiehi
XFILLER_19_934 VPWR VGND sg13g2_decap_8
XFILLER_46_775 VPWR VGND sg13g2_decap_8
XFILLER_45_252 VPWR VGND sg13g2_decap_4
XFILLER_33_403 VPWR VGND sg13g2_fill_2
XFILLER_33_447 VPWR VGND sg13g2_fill_1
XFILLER_33_469 VPWR VGND sg13g2_fill_1
XFILLER_9_131 VPWR VGND sg13g2_decap_4
XFILLER_13_171 VPWR VGND sg13g2_fill_1
X_3650_ net540 _0648_ mydesign.accum\[113\] _0663_ VPWR VGND sg13g2_nand3_1
X_3581_ _0606_ _0604_ _0605_ VPWR VGND sg13g2_nand2_1
X_5320_ net638 VPWR _2139_ VGND net520 net450 sg13g2_o21ai_1
X_5251_ _2009_ mydesign.pe_weights\[31\] _2081_ VPWR VGND sg13g2_nor2b_1
X_4202_ _1158_ _2572_ _1157_ VPWR VGND sg13g2_xnor2_1
X_5182_ net497 mydesign.inputs\[3\]\[7\] _2017_ VPWR VGND sg13g2_nor2_1
X_4133_ _1093_ _1092_ _1091_ VPWR VGND sg13g2_nand2b_1
X_4064_ net464 VPWR _1036_ VGND net566 net944 sg13g2_o21ai_1
XFILLER_28_208 VPWR VGND sg13g2_fill_1
XFILLER_24_425 VPWR VGND sg13g2_fill_1
XFILLER_25_959 VPWR VGND sg13g2_decap_8
X_4966_ _1799_ _1820_ _1821_ VPWR VGND sg13g2_nor2b_1
X_4897_ _2591_ _2648_ _2657_ _1767_ VPWR VGND sg13g2_nor3_2
XFILLER_20_631 VPWR VGND sg13g2_fill_1
XFILLER_22_15 VPWR VGND sg13g2_decap_4
X_3917_ VGND VPWR _0892_ _0901_ _0904_ _0900_ sg13g2_a21oi_1
X_3848_ mydesign.pe_inputs\[56\] VPWR _0839_ VGND _0800_ _0803_ sg13g2_o21ai_1
XFILLER_22_37 VPWR VGND sg13g2_decap_8
X_3779_ net622 VPWR _0778_ VGND mydesign.pe_inputs\[55\] net435 sg13g2_o21ai_1
X_5518_ VGND VPWR mydesign.pe_inputs\[11\] net525 _2319_ mydesign.accum\[13\] sg13g2_a21oi_1
XFILLER_0_8 VPWR VGND sg13g2_decap_4
X_5449_ _2252_ VPWR _2254_ VGND _2250_ _2251_ sg13g2_o21ai_1
XFILLER_43_701 VPWR VGND sg13g2_decap_4
XFILLER_27_241 VPWR VGND sg13g2_fill_1
XFILLER_28_764 VPWR VGND sg13g2_fill_1
XFILLER_43_767 VPWR VGND sg13g2_decap_8
XFILLER_42_222 VPWR VGND sg13g2_decap_8
XFILLER_24_981 VPWR VGND sg13g2_decap_8
XFILLER_31_929 VPWR VGND sg13g2_decap_8
XFILLER_11_642 VPWR VGND sg13g2_fill_1
XFILLER_6_112 VPWR VGND sg13g2_fill_2
XFILLER_3_830 VPWR VGND sg13g2_decap_8
XFILLER_3_863 VPWR VGND sg13g2_fill_1
XFILLER_3_885 VPWR VGND sg13g2_decap_4
XFILLER_19_764 VPWR VGND sg13g2_fill_1
XFILLER_46_572 VPWR VGND sg13g2_fill_2
XFILLER_19_786 VPWR VGND sg13g2_fill_1
XFILLER_33_211 VPWR VGND sg13g2_decap_4
XFILLER_22_918 VPWR VGND sg13g2_fill_1
XFILLER_33_233 VPWR VGND sg13g2_fill_1
XFILLER_33_244 VPWR VGND sg13g2_fill_1
X_4820_ _1684_ _1698_ _1699_ VPWR VGND sg13g2_and2_1
XFILLER_34_745 VPWR VGND sg13g2_fill_2
XFILLER_34_778 VPWR VGND sg13g2_decap_8
X_4751_ VGND VPWR _1630_ _1639_ _1642_ _1638_ sg13g2_a21oi_1
X_4682_ net535 VPWR _1577_ VGND _1517_ _1520_ sg13g2_o21ai_1
XFILLER_30_962 VPWR VGND sg13g2_decap_8
X_3702_ _0712_ _0694_ _0692_ VPWR VGND sg13g2_nand2b_1
X_3633_ VGND VPWR _2566_ net492 _0101_ _0649_ sg13g2_a21oi_1
X_3564_ _0590_ _0578_ _0588_ VPWR VGND sg13g2_xnor2_1
X_5303_ VGND VPWR net567 _2128_ _0291_ _2129_ sg13g2_a21oi_1
X_3495_ _2586_ _0525_ _0526_ VPWR VGND sg13g2_and2_1
X_5234_ _2063_ _2064_ _2040_ _2065_ VPWR VGND sg13g2_nand3_1
X_5165_ _2003_ net541 mydesign.inputs\[3\]\[0\] net496 VPWR VGND sg13g2_and3_1
X_4116_ VGND VPWR mydesign.accum\[88\] _1067_ _1077_ _1075_ sg13g2_a21oi_1
X_5096_ _1938_ _1921_ _1939_ VPWR VGND sg13g2_nor2b_1
X_4047_ _1019_ _1007_ _1020_ VPWR VGND sg13g2_xor2_1
XFILLER_33_14 VPWR VGND sg13g2_decap_8
X_5998_ net102 VGND VPWR _0224_ mydesign.accum\[60\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_40_759 VPWR VGND sg13g2_fill_2
X_4949_ _1787_ _1803_ _1805_ VPWR VGND sg13g2_nor2_1
XFILLER_33_47 VPWR VGND sg13g2_fill_1
XFILLER_32_1006 VPWR VGND sg13g2_decap_8
XFILLER_21_995 VPWR VGND sg13g2_decap_8
XFILLER_4_649 VPWR VGND sg13g2_decap_4
XFILLER_4_627 VPWR VGND sg13g2_decap_4
XFILLER_0_866 VPWR VGND sg13g2_decap_8
XFILLER_48_804 VPWR VGND sg13g2_decap_8
XFILLER_16_734 VPWR VGND sg13g2_fill_2
XFILLER_28_583 VPWR VGND sg13g2_fill_1
XFILLER_15_288 VPWR VGND sg13g2_fill_2
X_6062__210 VPWR VGND net210 sg13g2_tiehi
XFILLER_8_911 VPWR VGND sg13g2_fill_2
XFILLER_8_966 VPWR VGND sg13g2_decap_8
XFILLER_12_984 VPWR VGND sg13g2_decap_8
X_3280_ net614 VPWR _2684_ VGND _2657_ _2683_ sg13g2_o21ai_1
XFILLER_39_826 VPWR VGND sg13g2_fill_1
XFILLER_24_4 VPWR VGND sg13g2_decap_4
X_5921_ net315 VGND VPWR _0147_ mydesign.accum\[103\] clknet_leaf_45_clk sg13g2_dfrbpq_2
XFILLER_34_553 VPWR VGND sg13g2_decap_4
X_5852_ net67 VGND VPWR net419 mydesign.inputs\[2\]\[14\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_5783_ net171 VGND VPWR net678 mydesign.weights\[2\]\[16\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_4803_ VGND VPWR net582 _1681_ _0238_ _1682_ sg13g2_a21oi_1
XFILLER_21_258 VPWR VGND sg13g2_decap_8
XFILLER_21_269 VPWR VGND sg13g2_fill_1
X_4734_ _1627_ _1606_ _1625_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_770 VPWR VGND sg13g2_decap_4
X_4665_ _1559_ _1558_ _1561_ VPWR VGND sg13g2_xor2_1
X_4596_ _1504_ _1502_ _1503_ VPWR VGND sg13g2_xnor2_1
X_3616_ VGND VPWR _2582_ net486 _0097_ _0636_ sg13g2_a21oi_1
X_3547_ _0553_ _0573_ _0551_ _0574_ VPWR VGND sg13g2_nand3_1
XFILLER_0_118 VPWR VGND sg13g2_fill_1
X_6074__136 VPWR VGND net136 sg13g2_tiehi
X_3478_ _0513_ _0499_ _0512_ net484 net1059 VPWR VGND sg13g2_a22oi_1
X_5217_ _2048_ _2031_ _2049_ VPWR VGND sg13g2_xor2_1
X_5148_ _1987_ _1986_ _1988_ VPWR VGND sg13g2_xor2_1
XFILLER_45_807 VPWR VGND sg13g2_decap_8
X_5079_ _1913_ VPWR _1922_ VGND _1906_ _1914_ sg13g2_o21ai_1
XFILLER_38_881 VPWR VGND sg13g2_decap_8
XFILLER_12_225 VPWR VGND sg13g2_fill_1
XFILLER_25_597 VPWR VGND sg13g2_fill_1
XFILLER_48_601 VPWR VGND sg13g2_decap_8
XFILLER_48_678 VPWR VGND sg13g2_decap_8
XFILLER_29_892 VPWR VGND sg13g2_decap_8
XFILLER_16_520 VPWR VGND sg13g2_decap_8
XFILLER_44_862 VPWR VGND sg13g2_decap_8
XFILLER_43_361 VPWR VGND sg13g2_fill_1
XFILLER_31_501 VPWR VGND sg13g2_fill_1
XFILLER_43_394 VPWR VGND sg13g2_fill_2
XFILLER_7_284 VPWR VGND sg13g2_fill_2
Xhold207 mydesign.accum\[38\] VPWR VGND net826 sg13g2_dlygate4sd3_1
X_4450_ _1373_ _1372_ _1375_ VPWR VGND sg13g2_xor2_1
Xhold229 _0142_ VPWR VGND net848 sg13g2_dlygate4sd3_1
XFILLER_7_295 VPWR VGND sg13g2_fill_1
X_3401_ VGND VPWR net504 _0446_ _0448_ _0447_ sg13g2_a21oi_1
X_4381_ _1309_ mydesign.pe_weights\[53\] mydesign.pe_inputs\[41\] VPWR VGND sg13g2_nand2_1
Xhold218 mydesign.accum\[31\] VPWR VGND net837 sg13g2_dlygate4sd3_1
X_3332_ VGND VPWR _0388_ _0387_ net548 sg13g2_or2_1
X_6120_ net76 VGND VPWR _0346_ mydesign.weights\[1\]\[10\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_6051_ net254 VGND VPWR _0277_ mydesign.accum\[37\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3263_ VGND VPWR _2520_ _2673_ _0029_ _2674_ sg13g2_a21oi_1
X_5002_ net531 mydesign.pe_inputs\[26\] mydesign.accum\[45\] _1855_ VPWR VGND sg13g2_nand3_1
X_3194_ net728 _2623_ net620 _2628_ VPWR VGND sg13g2_nand3_1
XFILLER_15_0 VPWR VGND sg13g2_fill_2
X_5862__49 VPWR VGND net49 sg13g2_tiehi
X_6009__54 VPWR VGND net54 sg13g2_tiehi
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
X_5904_ net345 VGND VPWR _0130_ mydesign.accum\[110\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_35_862 VPWR VGND sg13g2_fill_1
XFILLER_35_873 VPWR VGND sg13g2_decap_8
X_5835_ net99 VGND VPWR _0061_ mydesign.compute_en clknet_leaf_47_clk sg13g2_dfrbpq_1
XFILLER_14_49 VPWR VGND sg13g2_fill_2
X_5766_ _2512_ net699 _2511_ VPWR VGND sg13g2_nand2_1
X_5697_ _2475_ VPWR _0339_ VGND net504 _2474_ sg13g2_o21ai_1
X_4717_ _1611_ _1593_ _1610_ VPWR VGND sg13g2_xnor2_1
X_4648_ mydesign.pe_weights\[45\] _1521_ mydesign.accum\[57\] _1545_ VPWR VGND sg13g2_nand3_1
X_4579_ _1466_ VPWR _1488_ VGND _1459_ _1467_ sg13g2_o21ai_1
XFILLER_39_24 VPWR VGND sg13g2_fill_2
XFILLER_39_13 VPWR VGND sg13g2_decap_8
X_5917__323 VPWR VGND net323 sg13g2_tiehi
XFILLER_17_328 VPWR VGND sg13g2_decap_8
XFILLER_44_114 VPWR VGND sg13g2_fill_1
XFILLER_26_851 VPWR VGND sg13g2_fill_2
X_5989__170 VPWR VGND net170 sg13g2_tiehi
XFILLER_40_320 VPWR VGND sg13g2_fill_2
XFILLER_26_895 VPWR VGND sg13g2_decap_4
XFILLER_13_578 VPWR VGND sg13g2_decap_4
X_6024__366 VPWR VGND net366 sg13g2_tiehi
XFILLER_5_700 VPWR VGND sg13g2_fill_1
X_6100__276 VPWR VGND net276 sg13g2_tiehi
XFILLER_20_92 VPWR VGND sg13g2_fill_2
XFILLER_1_950 VPWR VGND sg13g2_decap_8
XFILLER_49_965 VPWR VGND sg13g2_decap_8
Xhold90 mydesign.inputs\[3\]\[0\] VPWR VGND net709 sg13g2_dlygate4sd3_1
XFILLER_36_604 VPWR VGND sg13g2_decap_8
XFILLER_36_648 VPWR VGND sg13g2_fill_2
X_3950_ _0929_ net547 mydesign.weights\[3\]\[7\] VPWR VGND sg13g2_nand2_1
X_5968__221 VPWR VGND net221 sg13g2_tiehi
X_3881_ _0869_ _0870_ _0871_ VPWR VGND sg13g2_nor2b_1
X_5620_ _2410_ mydesign.pe_inputs\[6\] mydesign.pe_weights\[18\] VPWR VGND sg13g2_nand2_1
XFILLER_31_386 VPWR VGND sg13g2_fill_2
XFILLER_32_887 VPWR VGND sg13g2_decap_8
X_5551_ _2350_ mydesign.accum\[15\] _2349_ VPWR VGND sg13g2_xnor2_1
X_4502_ _1415_ mydesign.pe_weights\[48\] mydesign.pe_inputs\[37\] VPWR VGND sg13g2_nand2_1
X_5482_ _2283_ _2262_ _2285_ VPWR VGND sg13g2_xor2_1
X_4433_ _1357_ _1356_ _1359_ VPWR VGND sg13g2_xor2_1
Xfanout506 net507 net506 VPWR VGND sg13g2_buf_8
X_4364_ net637 VPWR _1295_ VGND net538 net493 sg13g2_o21ai_1
X_4295_ _1237_ _1231_ _1236_ VPWR VGND sg13g2_nand2_1
Xfanout539 net1096 net539 VPWR VGND sg13g2_buf_8
X_6103_ net252 VGND VPWR _0329_ mydesign.accum\[5\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3315_ _2603_ net431 _0376_ VPWR VGND sg13g2_nor2_1
Xfanout517 net518 net517 VPWR VGND sg13g2_buf_8
Xfanout528 net1022 net528 VPWR VGND sg13g2_buf_8
XFILLER_6_1021 VPWR VGND sg13g2_decap_8
X_6034_ net322 VGND VPWR net665 mydesign.accum\[40\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3246_ VGND VPWR _2662_ _2666_ _2665_ _2664_ sg13g2_a21oi_2
X_3177_ _2613_ VPWR _0003_ VGND net432 _2614_ sg13g2_o21ai_1
XFILLER_27_604 VPWR VGND sg13g2_fill_2
XFILLER_27_615 VPWR VGND sg13g2_decap_8
XFILLER_27_637 VPWR VGND sg13g2_decap_8
XFILLER_42_607 VPWR VGND sg13g2_fill_2
X_5818_ net124 VGND VPWR _0044_ mydesign.inputs\[1\]\[23\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_10_537 VPWR VGND sg13g2_fill_1
X_5749_ _2504_ net751 _2500_ VPWR VGND sg13g2_nand2_1
X_5882__385 VPWR VGND net385 sg13g2_tiehi
XFILLER_2_769 VPWR VGND sg13g2_fill_2
XFILLER_49_239 VPWR VGND sg13g2_decap_8
XFILLER_49_217 VPWR VGND sg13g2_decap_4
XFILLER_18_615 VPWR VGND sg13g2_decap_8
XFILLER_46_957 VPWR VGND sg13g2_decap_8
XFILLER_45_489 VPWR VGND sg13g2_fill_1
XFILLER_14_865 VPWR VGND sg13g2_fill_2
XFILLER_32_139 VPWR VGND sg13g2_fill_1
XFILLER_9_368 VPWR VGND sg13g2_fill_2
XFILLER_9_379 VPWR VGND sg13g2_fill_1
XFILLER_12_1026 VPWR VGND sg13g2_fill_2
X_5820__122 VPWR VGND net122 sg13g2_tiehi
X_3100_ VPWR _2541_ net789 VGND sg13g2_inv_1
X_4080_ _1049_ net544 net554 mydesign.inputs\[1\]\[13\] VPWR VGND sg13g2_and3_1
XFILLER_49_762 VPWR VGND sg13g2_decap_8
XFILLER_37_924 VPWR VGND sg13g2_decap_8
XFILLER_36_467 VPWR VGND sg13g2_decap_4
X_4982_ net531 mydesign.pe_inputs\[25\] mydesign.accum\[44\] _1836_ VPWR VGND sg13g2_nand3_1
X_3933_ net628 VPWR _0915_ VGND net1091 net433 sg13g2_o21ai_1
X_3864_ VGND VPWR net572 _0853_ _0127_ _0854_ sg13g2_a21oi_1
X_5603_ VGND VPWR net519 net523 _2394_ mydesign.accum\[3\] sg13g2_a21oi_1
X_3795_ _0791_ net551 mydesign.weights\[2\]\[6\] VPWR VGND sg13g2_nand2b_1
X_5534_ net520 mydesign.pe_weights\[23\] mydesign.accum\[14\] _2334_ VPWR VGND sg13g2_nand3_1
X_5465_ _2266_ _2250_ _2269_ VPWR VGND sg13g2_xor2_1
X_4416_ net474 VPWR _1343_ VGND net575 net868 sg13g2_o21ai_1
X_5396_ mydesign.pe_inputs\[14\] net527 mydesign.accum\[21\] _2209_ VPWR VGND sg13g2_nand3_1
X_4347_ _1285_ _1282_ _1286_ VPWR VGND sg13g2_xor2_1
X_4278_ _1219_ _1212_ _1221_ VPWR VGND sg13g2_xor2_1
X_6017_ net398 VGND VPWR _0243_ mydesign.accum\[55\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_39_261 VPWR VGND sg13g2_decap_4
X_3229_ _2652_ net413 _2650_ VPWR VGND sg13g2_nand2_1
XFILLER_28_935 VPWR VGND sg13g2_decap_8
XFILLER_43_949 VPWR VGND sg13g2_decap_8
XFILLER_2_533 VPWR VGND sg13g2_decap_8
XFILLER_2_500 VPWR VGND sg13g2_fill_1
XFILLER_2_544 VPWR VGND sg13g2_decap_4
Xhold390 mydesign.accum\[107\] VPWR VGND net1009 sg13g2_dlygate4sd3_1
XFILLER_46_754 VPWR VGND sg13g2_decap_8
XFILLER_27_990 VPWR VGND sg13g2_decap_8
XFILLER_33_415 VPWR VGND sg13g2_decap_8
XFILLER_34_949 VPWR VGND sg13g2_decap_8
XFILLER_42_982 VPWR VGND sg13g2_decap_8
XFILLER_14_684 VPWR VGND sg13g2_decap_8
X_3580_ _0582_ VPWR _0605_ VGND _0581_ _0584_ sg13g2_o21ai_1
XFILLER_10_890 VPWR VGND sg13g2_fill_1
XFILLER_6_861 VPWR VGND sg13g2_fill_1
X_5250_ _2080_ mydesign.pe_weights\[30\] _2015_ VPWR VGND sg13g2_nand2_1
X_4201_ _1157_ mydesign.pe_weights\[63\] _1061_ VPWR VGND sg13g2_nand2_1
X_6037__310 VPWR VGND net310 sg13g2_tiehi
X_5181_ VGND VPWR _2526_ net494 _0282_ _2016_ sg13g2_a21oi_1
X_4132_ VGND VPWR _1092_ _1090_ _1074_ sg13g2_or2_1
XFILLER_3_62 VPWR VGND sg13g2_fill_1
X_4063_ _1035_ _1023_ _1034_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_1013 VPWR VGND sg13g2_decap_8
XFILLER_25_927 VPWR VGND sg13g2_fill_2
XFILLER_25_938 VPWR VGND sg13g2_decap_8
X_4965_ _1819_ _1816_ _1820_ VPWR VGND sg13g2_xor2_1
XFILLER_11_109 VPWR VGND sg13g2_fill_2
X_3916_ VGND VPWR net570 _0902_ _0130_ _0903_ sg13g2_a21oi_1
X_4896_ _1766_ VPWR _0247_ VGND net597 _1761_ sg13g2_o21ai_1
XFILLER_32_492 VPWR VGND sg13g2_fill_2
X_3847_ _0838_ mydesign.pe_inputs\[57\] _0796_ VPWR VGND sg13g2_nand2_1
XFILLER_20_665 VPWR VGND sg13g2_decap_4
X_3778_ VGND VPWR _2581_ net435 _0118_ _0777_ sg13g2_a21oi_1
X_5517_ net520 net525 mydesign.accum\[13\] _2318_ VPWR VGND sg13g2_nand3_1
X_5448_ _2250_ _2251_ _2252_ _2253_ VPWR VGND sg13g2_nor3_1
X_5379_ _2193_ _2191_ _2192_ VPWR VGND sg13g2_nand2_1
XFILLER_47_529 VPWR VGND sg13g2_fill_1
XFILLER_27_253 VPWR VGND sg13g2_decap_8
XFILLER_16_949 VPWR VGND sg13g2_decap_8
XFILLER_27_275 VPWR VGND sg13g2_decap_8
XFILLER_43_746 VPWR VGND sg13g2_decap_8
XFILLER_15_459 VPWR VGND sg13g2_fill_2
XFILLER_31_908 VPWR VGND sg13g2_decap_8
XFILLER_24_960 VPWR VGND sg13g2_decap_8
XFILLER_10_120 VPWR VGND sg13g2_fill_1
XFILLER_6_135 VPWR VGND sg13g2_fill_1
XFILLER_6_102 VPWR VGND sg13g2_fill_1
XFILLER_10_186 VPWR VGND sg13g2_fill_2
XFILLER_6_157 VPWR VGND sg13g2_fill_1
XFILLER_26_8 VPWR VGND sg13g2_fill_1
XFILLER_19_721 VPWR VGND sg13g2_fill_1
XFILLER_34_724 VPWR VGND sg13g2_decap_4
XFILLER_33_278 VPWR VGND sg13g2_decap_4
X_4750_ VGND VPWR net567 _1640_ _0226_ _1641_ sg13g2_a21oi_1
XFILLER_15_993 VPWR VGND sg13g2_decap_8
XFILLER_30_941 VPWR VGND sg13g2_decap_8
X_3701_ _0711_ mydesign.pe_inputs\[63\] _0648_ VPWR VGND sg13g2_nand2_1
X_4681_ _1576_ mydesign.pe_weights\[46\] _1527_ VPWR VGND sg13g2_nand2_1
X_3632_ net631 VPWR _0649_ VGND net492 _0648_ sg13g2_o21ai_1
X_3563_ _0589_ _0578_ _0588_ VPWR VGND sg13g2_nand2_1
X_5302_ net470 VPWR _2129_ VGND net568 net837 sg13g2_o21ai_1
XFILLER_45_0 VPWR VGND sg13g2_decap_4
X_3494_ net556 mydesign.weights\[0\]\[27\] mydesign.weights\[0\]\[23\] mydesign.weights\[0\]\[19\]
+ mydesign.weights\[0\]\[15\] net545 _0525_ VPWR VGND sg13g2_mux4_1
X_5233_ _2062_ _2061_ _2055_ _2064_ VPWR VGND sg13g2_a21o_1
X_5164_ _2002_ net549 mydesign.inputs\[3\]\[12\] _0392_ VPWR VGND sg13g2_and3_1
X_4115_ _1076_ mydesign.accum\[88\] _1067_ _1075_ VPWR VGND sg13g2_and3_2
X_5095_ _1938_ _1922_ _1936_ VPWR VGND sg13g2_xnor2_1
X_4046_ _1019_ _0998_ _1018_ VPWR VGND sg13g2_xnor2_1
X_5997_ net106 VGND VPWR _0223_ mydesign.accum\[59\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_4948_ _1804_ _1787_ _1803_ VPWR VGND sg13g2_nand2_1
XFILLER_33_59 VPWR VGND sg13g2_decap_8
X_4879_ _1753_ _1754_ _0242_ VPWR VGND sg13g2_nor2_1
XFILLER_21_974 VPWR VGND sg13g2_decap_8
XFILLER_0_845 VPWR VGND sg13g2_decap_8
XFILLER_43_510 VPWR VGND sg13g2_fill_1
XFILLER_28_595 VPWR VGND sg13g2_fill_1
XFILLER_43_576 VPWR VGND sg13g2_fill_1
X_5927__303 VPWR VGND net303 sg13g2_tiehi
XFILLER_12_963 VPWR VGND sg13g2_decap_8
XFILLER_7_455 VPWR VGND sg13g2_decap_8
X_6103__252 VPWR VGND net252 sg13g2_tiehi
XFILLER_48_1014 VPWR VGND sg13g2_decap_8
X_5859__55 VPWR VGND net55 sg13g2_tiehi
X_5874__25 VPWR VGND net25 sg13g2_tiehi
XFILLER_38_359 VPWR VGND sg13g2_fill_2
X_6110__212 VPWR VGND net212 sg13g2_tiehi
XFILLER_0_41 VPWR VGND sg13g2_fill_2
XFILLER_0_1027 VPWR VGND sg13g2_fill_2
X_5920_ net317 VGND VPWR _0146_ mydesign.accum\[102\] clknet_leaf_45_clk sg13g2_dfrbpq_2
X_5851_ net68 VGND VPWR net426 mydesign.inputs\[2\]\[13\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_21_215 VPWR VGND sg13g2_decap_8
XFILLER_21_237 VPWR VGND sg13g2_fill_1
XFILLER_22_749 VPWR VGND sg13g2_decap_8
X_5782_ net172 VGND VPWR _0008_ mydesign.inputs\[0\]\[27\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_4802_ net479 VPWR _1682_ VGND net582 net900 sg13g2_o21ai_1
X_4733_ VGND VPWR _1626_ _1625_ _1606_ sg13g2_or2_1
X_4664_ _1558_ _1559_ _1560_ VPWR VGND sg13g2_nor2_1
X_5978__201 VPWR VGND net201 sg13g2_tiehi
X_4595_ _1503_ _1489_ _1486_ VPWR VGND sg13g2_nand2b_1
X_3615_ net630 VPWR _0636_ VGND mydesign.pe_inputs\[61\] net487 sg13g2_o21ai_1
X_3546_ _0573_ _0556_ _0571_ VPWR VGND sg13g2_xnor2_1
X_5216_ _2048_ _2047_ _2046_ VPWR VGND sg13g2_nand2b_1
X_3477_ _0511_ VPWR _0512_ VGND net544 _0510_ sg13g2_o21ai_1
X_5147_ VGND VPWR _1963_ _1971_ _1987_ _1970_ sg13g2_a21oi_1
XFILLER_29_315 VPWR VGND sg13g2_decap_8
X_5078_ _1917_ VPWR _1921_ VGND _1903_ _1918_ sg13g2_o21ai_1
XFILLER_28_59 VPWR VGND sg13g2_fill_2
X_4029_ VGND VPWR _0963_ _0983_ _1003_ _0982_ sg13g2_a21oi_1
XFILLER_44_69 VPWR VGND sg13g2_fill_2
XFILLER_21_782 VPWR VGND sg13g2_decap_4
XFILLER_5_915 VPWR VGND sg13g2_fill_1
XFILLER_4_425 VPWR VGND sg13g2_decap_4
XFILLER_0_664 VPWR VGND sg13g2_decap_4
XFILLER_48_657 VPWR VGND sg13g2_decap_8
XFILLER_44_841 VPWR VGND sg13g2_decap_8
XFILLER_16_510 VPWR VGND sg13g2_fill_1
XFILLER_43_384 VPWR VGND sg13g2_fill_1
XFILLER_31_524 VPWR VGND sg13g2_fill_2
Xhold208 mydesign.accum\[54\] VPWR VGND net827 sg13g2_dlygate4sd3_1
Xhold219 mydesign.pe_weights\[62\] VPWR VGND net838 sg13g2_dlygate4sd3_1
X_3400_ net458 VPWR _0447_ VGND net504 _0444_ sg13g2_o21ai_1
X_4380_ _1308_ mydesign.pe_weights\[52\] mydesign.pe_inputs\[42\] VPWR VGND sg13g2_nand2_1
X_3331_ VGND VPWR _2604_ _0387_ _2598_ net454 sg13g2_a21oi_2
XFILLER_39_602 VPWR VGND sg13g2_decap_8
X_6050_ net258 VGND VPWR _0276_ mydesign.accum\[36\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3262_ net617 VPWR _2674_ VGND net805 _2673_ sg13g2_o21ai_1
X_5001_ _1854_ mydesign.pe_weights\[38\] mydesign.pe_inputs\[27\] VPWR VGND sg13g2_nand2_1
X_3193_ _2626_ VPWR _0006_ VGND _2623_ net601 sg13g2_o21ai_1
XFILLER_38_101 VPWR VGND sg13g2_fill_1
XFILLER_39_668 VPWR VGND sg13g2_fill_2
XFILLER_22_1017 VPWR VGND sg13g2_decap_8
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
X_5903_ net347 VGND VPWR _0129_ mydesign.accum\[109\] clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_35_852 VPWR VGND sg13g2_fill_2
X_5834_ net101 VGND VPWR _0060_ mydesign.load_counter\[3\] clknet_leaf_1_clk sg13g2_dfrbpq_2
XFILLER_22_579 VPWR VGND sg13g2_fill_2
X_5765_ _2511_ net462 _0910_ VPWR VGND sg13g2_nand2_2
X_5696_ net504 VPWR _2475_ VGND _2466_ _2471_ sg13g2_o21ai_1
X_4716_ _1610_ _1607_ _1608_ VPWR VGND sg13g2_xnor2_1
X_4647_ VGND VPWR net686 _1543_ _0220_ _1544_ sg13g2_a21oi_1
X_4578_ _1485_ _1484_ _1487_ VPWR VGND sg13g2_xor2_1
X_5798__152 VPWR VGND net152 sg13g2_tiehi
X_3529_ _0556_ _0547_ _0549_ VPWR VGND sg13g2_nand2_1
XFILLER_29_189 VPWR VGND sg13g2_decap_8
XFILLER_41_888 VPWR VGND sg13g2_decap_8
XFILLER_4_266 VPWR VGND sg13g2_fill_2
XFILLER_45_1017 VPWR VGND sg13g2_decap_8
XFILLER_4_299 VPWR VGND sg13g2_decap_4
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_944 VPWR VGND sg13g2_decap_8
XFILLER_0_472 VPWR VGND sg13g2_decap_8
Xhold91 _0053_ VPWR VGND net710 sg13g2_dlygate4sd3_1
Xhold80 mydesign.weights\[1\]\[20\] VPWR VGND net699 sg13g2_dlygate4sd3_1
XFILLER_36_616 VPWR VGND sg13g2_fill_1
XFILLER_29_690 VPWR VGND sg13g2_fill_1
XFILLER_35_115 VPWR VGND sg13g2_fill_1
X_3880_ _0847_ VPWR _0870_ VGND _0836_ _0848_ sg13g2_o21ai_1
X_5550_ _2334_ VPWR _2349_ VGND _2333_ _2337_ sg13g2_o21ai_1
XFILLER_8_572 VPWR VGND sg13g2_fill_1
XFILLER_8_561 VPWR VGND sg13g2_decap_8
X_4501_ VGND VPWR mydesign.pe_weights\[49\] net532 _1414_ mydesign.accum\[65\] sg13g2_a21oi_1
X_5481_ _2262_ _2283_ _2284_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_594 VPWR VGND sg13g2_fill_1
X_4432_ _1358_ _1356_ _1357_ VPWR VGND sg13g2_nand2_1
X_4363_ VGND VPWR _2557_ net441 _0186_ _1294_ sg13g2_a21oi_1
X_4294_ _1235_ _1232_ _1236_ VPWR VGND sg13g2_xor2_1
X_6102_ net260 VGND VPWR _0328_ mydesign.accum\[4\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3314_ net6 _2599_ net499 _2698_ VPWR VGND sg13g2_nand3_1
Xfanout507 net510 net507 VPWR VGND sg13g2_buf_8
Xfanout518 net1105 net518 VPWR VGND sg13g2_buf_8
Xfanout529 net1094 net529 VPWR VGND sg13g2_buf_8
XFILLER_39_410 VPWR VGND sg13g2_decap_4
XFILLER_6_1000 VPWR VGND sg13g2_decap_8
X_3245_ _2588_ VPWR _2665_ VGND net596 mydesign.load_counter\[0\] sg13g2_o21ai_1
X_6033_ net326 VGND VPWR net1026 mydesign.pe_weights\[23\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_3176_ _2614_ net741 net616 VPWR VGND sg13g2_nand2_1
X_5843__83 VPWR VGND net83 sg13g2_tiehi
XFILLER_26_137 VPWR VGND sg13g2_fill_2
XFILLER_34_170 VPWR VGND sg13g2_fill_1
X_5817_ net125 VGND VPWR _0043_ mydesign.inputs\[1\]\[22\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_22_354 VPWR VGND sg13g2_decap_8
XFILLER_22_376 VPWR VGND sg13g2_decap_8
XFILLER_41_26 VPWR VGND sg13g2_fill_1
X_5748_ _2503_ VPWR _0362_ VGND _1773_ _2500_ sg13g2_o21ai_1
X_5679_ _2463_ VPWR _0333_ VGND net602 _2461_ sg13g2_o21ai_1
X_6093__332 VPWR VGND net332 sg13g2_tiehi
XFILLER_49_207 VPWR VGND sg13g2_fill_1
XFILLER_46_936 VPWR VGND sg13g2_decap_8
XFILLER_45_468 VPWR VGND sg13g2_fill_2
XFILLER_41_630 VPWR VGND sg13g2_fill_2
XFILLER_13_343 VPWR VGND sg13g2_fill_1
XFILLER_15_93 VPWR VGND sg13g2_decap_8
XFILLER_40_195 VPWR VGND sg13g2_decap_8
XFILLER_12_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_49_741 VPWR VGND sg13g2_decap_8
XFILLER_37_903 VPWR VGND sg13g2_decap_8
X_5935__287 VPWR VGND net287 sg13g2_tiehi
X_4981_ _1835_ mydesign.pe_weights\[38\] mydesign.pe_inputs\[26\] VPWR VGND sg13g2_nand2_1
XFILLER_23_118 VPWR VGND sg13g2_fill_2
X_3932_ VPWR VGND net985 _0913_ _0395_ net725 _0914_ net454 sg13g2_a221oi_1
Xclkbuf_leaf_43_clk clknet_3_4__leaf_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
XFILLER_17_693 VPWR VGND sg13g2_decap_8
XFILLER_32_630 VPWR VGND sg13g2_decap_4
X_3863_ net465 VPWR _0854_ VGND net572 net1009 sg13g2_o21ai_1
X_5788__162 VPWR VGND net162 sg13g2_tiehi
X_5602_ mydesign.pe_inputs\[7\] net523 mydesign.accum\[3\] _2393_ VPWR VGND sg13g2_nand3_1
X_3794_ VGND VPWR _2558_ net491 _0121_ _0790_ sg13g2_a21oi_1
X_5533_ VGND VPWR net520 mydesign.pe_weights\[23\] _2333_ mydesign.accum\[14\] sg13g2_a21oi_1
X_5464_ _2250_ _2266_ _2268_ VPWR VGND sg13g2_nor2_1
X_5395_ _2208_ mydesign.pe_inputs\[15\] mydesign.pe_weights\[26\] VPWR VGND sg13g2_nand2_1
X_4415_ _1340_ _1323_ _1342_ VPWR VGND sg13g2_xor2_1
X_4346_ _1285_ _1273_ _1284_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_1012 VPWR VGND sg13g2_decap_8
X_5795__155 VPWR VGND net155 sg13g2_tiehi
X_4277_ _1212_ _1219_ _1220_ VPWR VGND sg13g2_nor2_1
X_6016_ net26 VGND VPWR _0242_ mydesign.accum\[54\] clknet_leaf_26_clk sg13g2_dfrbpq_2
XFILLER_39_240 VPWR VGND sg13g2_fill_1
X_3228_ _2651_ VPWR _0017_ VGND net604 _2649_ sg13g2_o21ai_1
XFILLER_39_295 VPWR VGND sg13g2_decap_4
X_3159_ VGND VPWR _2600_ net5 net610 sg13g2_or2_1
XFILLER_43_928 VPWR VGND sg13g2_decap_8
XFILLER_14_118 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_34_clk clknet_3_5__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
XFILLER_11_825 VPWR VGND sg13g2_decap_4
XFILLER_23_663 VPWR VGND sg13g2_fill_1
X_5986__185 VPWR VGND net185 sg13g2_tiehi
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
Xhold380 mydesign.accum\[93\] VPWR VGND net999 sg13g2_dlygate4sd3_1
Xhold391 mydesign.accum\[106\] VPWR VGND net1010 sg13g2_dlygate4sd3_1
XFILLER_46_733 VPWR VGND sg13g2_decap_8
XFILLER_18_413 VPWR VGND sg13g2_fill_1
XFILLER_18_446 VPWR VGND sg13g2_decap_4
XFILLER_19_969 VPWR VGND sg13g2_decap_8
XFILLER_33_405 VPWR VGND sg13g2_fill_1
XFILLER_34_928 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_25_clk clknet_3_6__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_33_438 VPWR VGND sg13g2_decap_4
XFILLER_42_961 VPWR VGND sg13g2_decap_8
X_4200_ _1144_ VPWR _1156_ VGND _2573_ _1142_ sg13g2_o21ai_1
X_5180_ net625 VPWR _2016_ VGND net487 _2015_ sg13g2_o21ai_1
X_4131_ _1074_ _1090_ _1091_ VPWR VGND sg13g2_and2_1
X_4062_ _1034_ _1017_ _1031_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_744 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_16_clk clknet_3_2__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_4964_ _1819_ _1817_ _1818_ VPWR VGND sg13g2_nand2_1
XFILLER_20_600 VPWR VGND sg13g2_decap_4
X_3915_ net470 VPWR _0903_ VGND net570 net998 sg13g2_o21ai_1
X_4895_ _1766_ net648 _1762_ VPWR VGND sg13g2_nand2_1
XFILLER_33_994 VPWR VGND sg13g2_decap_8
X_3846_ _0837_ mydesign.pe_inputs\[58\] _0789_ VPWR VGND sg13g2_nand2_1
XFILLER_20_655 VPWR VGND sg13g2_fill_1
X_3777_ net627 VPWR _0777_ VGND net1036 net433 sg13g2_o21ai_1
X_5516_ _2317_ mydesign.accum\[13\] net520 net525 VPWR VGND sg13g2_and3_1
X_5447_ _2252_ mydesign.pe_inputs\[9\] mydesign.pe_weights\[20\] VPWR VGND sg13g2_nand2_1
X_5378_ net527 mydesign.pe_inputs\[13\] mydesign.accum\[20\] _2192_ VPWR VGND sg13g2_a21o_1
X_4329_ _1269_ _1268_ _1267_ VPWR VGND sg13g2_nand2b_1
XFILLER_43_725 VPWR VGND sg13g2_decap_8
XFILLER_27_265 VPWR VGND sg13g2_fill_2
X_5810__133 VPWR VGND net133 sg13g2_tiehi
XFILLER_10_143 VPWR VGND sg13g2_decap_4
XFILLER_6_114 VPWR VGND sg13g2_fill_1
XFILLER_5_0 VPWR VGND sg13g2_fill_1
X_5895__363 VPWR VGND net363 sg13g2_tiehi
XFILLER_38_508 VPWR VGND sg13g2_decap_8
XFILLER_34_747 VPWR VGND sg13g2_fill_1
XFILLER_15_972 VPWR VGND sg13g2_decap_8
XFILLER_42_791 VPWR VGND sg13g2_decap_8
XFILLER_30_920 VPWR VGND sg13g2_decap_8
X_3700_ _0696_ _0698_ _0710_ VPWR VGND sg13g2_nor2b_1
X_4680_ VPWR _1575_ _1574_ VGND sg13g2_inv_1
XFILLER_30_997 VPWR VGND sg13g2_decap_8
X_3631_ _0639_ net774 _0647_ _0648_ VPWR VGND sg13g2_a21o_2
X_3562_ _0587_ _0579_ _0588_ VPWR VGND sg13g2_xor2_1
X_5301_ _2127_ _2124_ _2128_ VPWR VGND sg13g2_xor2_1
X_3493_ VGND VPWR _2576_ net485 _0086_ _0524_ sg13g2_a21oi_1
Xclkbuf_leaf_5_clk clknet_3_1__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_5232_ _2061_ _2062_ _2055_ _2063_ VPWR VGND sg13g2_nand3_1
X_5163_ _0397_ _1999_ _2000_ _2001_ VPWR VGND sg13g2_nor3_1
XFILLER_25_1015 VPWR VGND sg13g2_decap_8
XFILLER_38_0 VPWR VGND sg13g2_decap_4
X_4114_ _1073_ _1072_ _1075_ VPWR VGND sg13g2_xor2_1
X_5094_ _1922_ _1936_ _1937_ VPWR VGND sg13g2_and2_1
X_5792__158 VPWR VGND net158 sg13g2_tiehi
XFILLER_49_390 VPWR VGND sg13g2_decap_8
X_4045_ _1018_ _1008_ _1016_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_585 VPWR VGND sg13g2_fill_2
X_5996_ net110 VGND VPWR _0222_ mydesign.accum\[58\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_4947_ _1801_ _1798_ _1803_ VPWR VGND sg13g2_xor2_1
XFILLER_33_780 VPWR VGND sg13g2_fill_1
X_4878_ net482 VPWR _1754_ VGND net582 net827 sg13g2_o21ai_1
XFILLER_20_441 VPWR VGND sg13g2_decap_4
XFILLER_21_953 VPWR VGND sg13g2_decap_8
X_3829_ _0819_ mydesign.accum\[106\] _0821_ VPWR VGND sg13g2_xor2_1
XFILLER_0_824 VPWR VGND sg13g2_decap_8
XFILLER_48_839 VPWR VGND sg13g2_decap_8
XFILLER_47_349 VPWR VGND sg13g2_decap_4
XFILLER_15_213 VPWR VGND sg13g2_fill_2
XFILLER_16_747 VPWR VGND sg13g2_fill_1
XFILLER_31_706 VPWR VGND sg13g2_fill_1
XFILLER_8_913 VPWR VGND sg13g2_fill_1
X_6027__354 VPWR VGND net354 sg13g2_tiehi
XFILLER_12_942 VPWR VGND sg13g2_decap_8
XFILLER_8_935 VPWR VGND sg13g2_fill_2
XFILLER_23_82 VPWR VGND sg13g2_fill_1
XFILLER_19_541 VPWR VGND sg13g2_decap_8
XFILLER_0_1006 VPWR VGND sg13g2_decap_8
XFILLER_19_552 VPWR VGND sg13g2_fill_2
XFILLER_47_894 VPWR VGND sg13g2_decap_8
X_5850_ net69 VGND VPWR net415 mydesign.inputs\[2\]\[12\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_5781_ net173 VGND VPWR _0007_ mydesign.inputs\[0\]\[26\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_4801_ _1681_ _1665_ _1680_ VPWR VGND sg13g2_xnor2_1
X_4732_ _1625_ _1623_ _1624_ VPWR VGND sg13g2_nand2_1
X_4663_ _1559_ mydesign.pe_weights\[45\] _1527_ VPWR VGND sg13g2_nand2_1
X_3614_ VGND VPWR _2583_ net486 _0096_ _0635_ sg13g2_a21oi_1
X_4594_ _1502_ _1501_ _1500_ VPWR VGND sg13g2_nand2b_1
X_3545_ _0572_ _0556_ _0571_ VPWR VGND sg13g2_nand2_1
X_3476_ _0511_ _0394_ mydesign.inputs\[0\]\[15\] net495 mydesign.inputs\[0\]\[19\]
+ VPWR VGND sg13g2_a22oi_1
X_5215_ VGND VPWR _2047_ _2045_ _2029_ sg13g2_or2_1
X_5146_ _1986_ _1985_ _1984_ VPWR VGND sg13g2_nand2b_1
X_5077_ VGND VPWR net584 _1919_ _0274_ _1920_ sg13g2_a21oi_1
XFILLER_44_308 VPWR VGND sg13g2_fill_2
X_4028_ _1000_ _0999_ _1002_ VPWR VGND sg13g2_xor2_1
X_5979_ net199 VGND VPWR net908 mydesign.accum\[65\] clknet_leaf_39_clk sg13g2_dfrbpq_2
XFILLER_21_794 VPWR VGND sg13g2_fill_1
XFILLER_0_643 VPWR VGND sg13g2_decap_8
XFILLER_48_636 VPWR VGND sg13g2_decap_8
XFILLER_0_687 VPWR VGND sg13g2_decap_8
XFILLER_0_698 VPWR VGND sg13g2_fill_2
XFILLER_47_146 VPWR VGND sg13g2_decap_8
XFILLER_44_820 VPWR VGND sg13g2_decap_8
XFILLER_44_897 VPWR VGND sg13g2_decap_8
XFILLER_16_577 VPWR VGND sg13g2_fill_2
XFILLER_43_396 VPWR VGND sg13g2_fill_1
XFILLER_34_70 VPWR VGND sg13g2_fill_1
XFILLER_15_1014 VPWR VGND sg13g2_decap_8
Xhold209 mydesign.pe_weights\[33\] VPWR VGND net828 sg13g2_dlygate4sd3_1
XFILLER_7_286 VPWR VGND sg13g2_fill_1
X_3330_ net607 _0386_ _0061_ VPWR VGND sg13g2_nor2_1
X_3261_ _2591_ _2671_ _2673_ VPWR VGND sg13g2_nor2_2
X_5000_ _1852_ _1853_ _0264_ VPWR VGND sg13g2_nor2_1
X_3192_ _2627_ net2 net620 VPWR VGND sg13g2_nand2_2
XFILLER_15_2 VPWR VGND sg13g2_fill_1
XFILLER_47_691 VPWR VGND sg13g2_decap_8
X_5902_ net349 VGND VPWR _0128_ mydesign.accum\[108\] clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_34_330 VPWR VGND sg13g2_fill_1
X_5833_ net103 VGND VPWR _0059_ mydesign.load_counter\[2\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5764_ net781 _2488_ _2510_ _0371_ VPWR VGND sg13g2_mux2_1
X_5945__267 VPWR VGND net267 sg13g2_tiehi
X_5695_ net457 _2467_ net512 _2474_ VPWR VGND sg13g2_nand3_1
XFILLER_30_591 VPWR VGND sg13g2_fill_2
X_4715_ VGND VPWR _1585_ _1587_ _1609_ _1607_ sg13g2_a21oi_1
X_4646_ net467 VPWR _1544_ VGND net686 _1543_ sg13g2_o21ai_1
X_4577_ _1484_ _1485_ _1486_ VPWR VGND sg13g2_and2_1
X_3528_ VGND VPWR net558 _0554_ _0090_ _0555_ sg13g2_a21oi_1
X_3459_ _0497_ VPWR _0079_ VGND net597 _0492_ sg13g2_o21ai_1
X_5129_ VGND VPWR _1945_ _1948_ _1970_ _1969_ sg13g2_a21oi_1
X_5861__51 VPWR VGND net51 sg13g2_tiehi
XFILLER_45_639 VPWR VGND sg13g2_decap_8
XFILLER_38_1014 VPWR VGND sg13g2_decap_8
XFILLER_26_853 VPWR VGND sg13g2_fill_1
XFILLER_13_503 VPWR VGND sg13g2_decap_8
XFILLER_41_867 VPWR VGND sg13g2_decap_8
XFILLER_40_322 VPWR VGND sg13g2_fill_1
XFILLER_9_529 VPWR VGND sg13g2_fill_2
XFILLER_5_713 VPWR VGND sg13g2_fill_2
X_5996__110 VPWR VGND net110 sg13g2_tiehi
XFILLER_4_234 VPWR VGND sg13g2_fill_2
XFILLER_49_923 VPWR VGND sg13g2_decap_8
XFILLER_1_985 VPWR VGND sg13g2_decap_8
XFILLER_48_466 VPWR VGND sg13g2_fill_2
Xhold70 _0124_ VPWR VGND net689 sg13g2_dlygate4sd3_1
Xhold92 mydesign.weights\[0\]\[26\] VPWR VGND net711 sg13g2_dlygate4sd3_1
Xhold81 mydesign.weights\[0\]\[21\] VPWR VGND net700 sg13g2_dlygate4sd3_1
XFILLER_17_820 VPWR VGND sg13g2_fill_1
XFILLER_17_853 VPWR VGND sg13g2_decap_4
XFILLER_44_694 VPWR VGND sg13g2_decap_8
XFILLER_43_160 VPWR VGND sg13g2_decap_8
XFILLER_32_801 VPWR VGND sg13g2_fill_2
XFILLER_32_812 VPWR VGND sg13g2_decap_8
X_4500_ _1413_ mydesign.accum\[65\] mydesign.pe_weights\[49\] net532 VPWR VGND sg13g2_and3_2
X_5480_ _2282_ _2279_ _2283_ VPWR VGND sg13g2_xor2_1
X_4431_ _1336_ VPWR _1357_ VGND _1325_ _1337_ sg13g2_o21ai_1
X_4362_ net636 VPWR _1294_ VGND net830 net441 sg13g2_o21ai_1
X_4293_ _1235_ _1233_ _1234_ VPWR VGND sg13g2_nand2_1
Xfanout519 mydesign.pe_inputs\[7\] net519 VPWR VGND sg13g2_buf_2
X_6101_ net268 VGND VPWR _0327_ mydesign.accum\[3\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3313_ _2697_ net499 net6 _2599_ VPWR VGND sg13g2_and3_1
Xfanout508 net509 net508 VPWR VGND sg13g2_buf_8
X_3244_ _2632_ _2663_ _2664_ VPWR VGND sg13g2_nor2_1
X_6032_ net330 VGND VPWR net831 mydesign.pe_weights\[22\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_3175_ _2613_ net3 net432 VPWR VGND sg13g2_nand2_1
XFILLER_27_628 VPWR VGND sg13g2_fill_1
XFILLER_23_834 VPWR VGND sg13g2_decap_8
XFILLER_35_672 VPWR VGND sg13g2_fill_2
XFILLER_35_683 VPWR VGND sg13g2_fill_1
X_5816_ net126 VGND VPWR _0042_ mydesign.inputs\[1\]\[21\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5747_ _2503_ net698 _2500_ VPWR VGND sg13g2_nand2_1
X_6127__392 VPWR VGND net392 sg13g2_tiehi
X_5678_ _2463_ net679 _2461_ VPWR VGND sg13g2_nand2_1
X_4629_ VGND VPWR net438 _1531_ _0214_ _1532_ sg13g2_a21oi_1
XFILLER_2_749 VPWR VGND sg13g2_fill_2
XFILLER_46_915 VPWR VGND sg13g2_decap_8
XFILLER_45_414 VPWR VGND sg13g2_decap_8
XFILLER_17_138 VPWR VGND sg13g2_fill_2
XFILLER_40_152 VPWR VGND sg13g2_fill_2
XFILLER_9_326 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_31_93 VPWR VGND sg13g2_fill_1
XFILLER_49_720 VPWR VGND sg13g2_decap_8
XFILLER_49_797 VPWR VGND sg13g2_decap_8
XFILLER_37_959 VPWR VGND sg13g2_decap_8
XFILLER_17_672 VPWR VGND sg13g2_decap_8
X_4980_ _1817_ VPWR _1834_ VGND _1816_ _1819_ sg13g2_o21ai_1
X_3931_ VGND VPWR net547 _2593_ _0913_ _0912_ sg13g2_a21oi_1
X_3862_ _0853_ _0834_ _0852_ VPWR VGND sg13g2_xnor2_1
X_5601_ _2392_ mydesign.accum\[3\] net519 net523 VPWR VGND sg13g2_and3_1
XFILLER_20_826 VPWR VGND sg13g2_decap_8
X_3793_ net629 VPWR _0790_ VGND net491 _0789_ sg13g2_o21ai_1
X_5532_ net463 _2332_ _0317_ VPWR VGND sg13g2_nor2_1
X_5463_ _2267_ _2250_ _2266_ VPWR VGND sg13g2_nand2_1
X_5394_ _2206_ _2207_ _0304_ VPWR VGND sg13g2_nor2_1
X_4414_ _1340_ _1323_ _1341_ VPWR VGND sg13g2_nor2b_1
X_4345_ _1284_ net865 _1283_ VPWR VGND sg13g2_xnor2_1
X_4276_ _1217_ _1196_ _1219_ VPWR VGND sg13g2_xor2_1
X_6015_ net30 VGND VPWR _0241_ mydesign.accum\[53\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_3227_ _2651_ net655 _2650_ VPWR VGND sg13g2_nand2_1
X_3158_ net610 net5 _2599_ VPWR VGND sg13g2_nor2_2
XFILLER_43_907 VPWR VGND sg13g2_decap_8
XFILLER_27_458 VPWR VGND sg13g2_fill_1
XFILLER_42_428 VPWR VGND sg13g2_fill_2
X_3089_ VPWR _2530_ net530 VGND sg13g2_inv_1
XFILLER_35_480 VPWR VGND sg13g2_fill_2
XFILLER_22_141 VPWR VGND sg13g2_fill_1
XFILLER_35_1006 VPWR VGND sg13g2_decap_8
XFILLER_23_697 VPWR VGND sg13g2_decap_8
XFILLER_2_513 VPWR VGND sg13g2_fill_2
Xhold370 mydesign.pe_weights\[57\] VPWR VGND net989 sg13g2_dlygate4sd3_1
XFILLER_7_4 VPWR VGND sg13g2_fill_2
XFILLER_2_557 VPWR VGND sg13g2_decap_8
Xhold381 mydesign.pe_inputs\[15\] VPWR VGND net1000 sg13g2_dlygate4sd3_1
Xhold392 _0126_ VPWR VGND net1011 sg13g2_dlygate4sd3_1
XFILLER_46_712 VPWR VGND sg13g2_decap_8
XFILLER_19_948 VPWR VGND sg13g2_decap_8
XFILLER_45_233 VPWR VGND sg13g2_decap_8
XFILLER_34_907 VPWR VGND sg13g2_decap_8
XFILLER_46_789 VPWR VGND sg13g2_decap_8
XFILLER_42_940 VPWR VGND sg13g2_decap_8
XFILLER_13_130 VPWR VGND sg13g2_fill_1
XFILLER_10_870 VPWR VGND sg13g2_decap_4
XFILLER_6_841 VPWR VGND sg13g2_fill_2
XFILLER_6_874 VPWR VGND sg13g2_fill_2
XFILLER_5_395 VPWR VGND sg13g2_decap_8
X_4130_ _1090_ _1080_ _1088_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_701 VPWR VGND sg13g2_fill_1
X_4061_ VPWR _1033_ _1032_ VGND sg13g2_inv_1
XFILLER_49_594 VPWR VGND sg13g2_decap_8
XFILLER_18_981 VPWR VGND sg13g2_decap_8
X_4963_ mydesign.pe_inputs\[24\] net531 mydesign.accum\[43\] _1818_ VPWR VGND sg13g2_a21o_1
X_3914_ _0902_ _0892_ _0901_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_450 VPWR VGND sg13g2_fill_1
XFILLER_33_973 VPWR VGND sg13g2_decap_8
X_4894_ _1765_ VPWR _0246_ VGND net599 _1761_ sg13g2_o21ai_1
X_3845_ _0836_ mydesign.pe_inputs\[59\] _0783_ VPWR VGND sg13g2_nand2_1
X_3776_ VGND VPWR _2582_ net433 _0117_ _0776_ sg13g2_a21oi_1
X_5515_ _2316_ mydesign.pe_inputs\[10\] mydesign.pe_weights\[23\] VPWR VGND sg13g2_nand2_1
X_5446_ VGND VPWR net521 mydesign.pe_weights\[21\] _2251_ mydesign.accum\[9\] sg13g2_a21oi_1
X_5377_ mydesign.pe_inputs\[13\] net527 mydesign.accum\[20\] _2191_ VPWR VGND sg13g2_nand3_1
X_4328_ net539 mydesign.pe_inputs\[47\] mydesign.accum\[86\] _1268_ VPWR VGND sg13g2_nand3_1
XFILLER_47_37 VPWR VGND sg13g2_fill_2
X_4259_ _1200_ _1184_ _1203_ VPWR VGND sg13g2_xor2_1
XFILLER_41_1021 VPWR VGND sg13g2_decap_8
XFILLER_27_222 VPWR VGND sg13g2_fill_2
XFILLER_42_236 VPWR VGND sg13g2_fill_1
XFILLER_27_299 VPWR VGND sg13g2_fill_1
XFILLER_23_450 VPWR VGND sg13g2_fill_2
XFILLER_24_995 VPWR VGND sg13g2_decap_8
XFILLER_11_634 VPWR VGND sg13g2_fill_1
XFILLER_10_188 VPWR VGND sg13g2_fill_1
XFILLER_2_332 VPWR VGND sg13g2_decap_4
XFILLER_2_354 VPWR VGND sg13g2_decap_8
XFILLER_2_387 VPWR VGND sg13g2_fill_1
XFILLER_18_211 VPWR VGND sg13g2_fill_1
XFILLER_15_951 VPWR VGND sg13g2_decap_8
XFILLER_18_1023 VPWR VGND sg13g2_decap_4
X_3630_ VGND VPWR _0645_ _0646_ _0647_ net542 sg13g2_a21oi_1
XFILLER_30_976 VPWR VGND sg13g2_decap_8
X_3561_ _0587_ _0580_ _0585_ VPWR VGND sg13g2_xnor2_1
X_5300_ _2127_ _2117_ _2126_ VPWR VGND sg13g2_xnor2_1
X_3492_ net624 VPWR _0524_ VGND net485 _0523_ sg13g2_o21ai_1
X_5231_ _2060_ _2059_ _2036_ _2062_ VPWR VGND sg13g2_a21o_1
X_5162_ net549 mydesign.inputs\[3\]\[8\] _2000_ VPWR VGND sg13g2_nor2_1
X_4113_ _1072_ _1073_ _1074_ VPWR VGND sg13g2_nor2_1
X_5093_ _1935_ _1923_ _1936_ VPWR VGND sg13g2_xor2_1
XFILLER_37_542 VPWR VGND sg13g2_fill_2
X_4044_ _1017_ _1008_ _1016_ VPWR VGND sg13g2_nand2_1
XFILLER_24_258 VPWR VGND sg13g2_fill_2
XFILLER_24_269 VPWR VGND sg13g2_fill_1
X_5995_ net114 VGND VPWR net819 mydesign.accum\[57\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_4946_ _1798_ _1801_ _1802_ VPWR VGND sg13g2_nor2_1
XFILLER_21_932 VPWR VGND sg13g2_decap_8
X_4877_ VGND VPWR _1751_ _1752_ _1753_ net502 sg13g2_a21oi_1
X_3828_ _0820_ mydesign.accum\[106\] _0819_ VPWR VGND sg13g2_nand2_1
X_3759_ _0766_ _0753_ _0765_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_129 VPWR VGND sg13g2_fill_1
X_5429_ _2240_ net978 _2226_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_803 VPWR VGND sg13g2_decap_8
XFILLER_48_818 VPWR VGND sg13g2_decap_8
X_5955__247 VPWR VGND net247 sg13g2_tiehi
XFILLER_12_921 VPWR VGND sg13g2_decap_8
XFILLER_12_998 VPWR VGND sg13g2_decap_8
XFILLER_7_468 VPWR VGND sg13g2_decap_4
XFILLER_3_663 VPWR VGND sg13g2_fill_1
XFILLER_3_641 VPWR VGND sg13g2_fill_1
XFILLER_47_873 VPWR VGND sg13g2_decap_8
XFILLER_0_43 VPWR VGND sg13g2_fill_1
XFILLER_19_575 VPWR VGND sg13g2_decap_4
XFILLER_34_523 VPWR VGND sg13g2_fill_2
X_4800_ _1680_ _1661_ _1678_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_228 VPWR VGND sg13g2_fill_1
X_5780_ net174 VGND VPWR _0006_ mydesign.inputs\[0\]\[25\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4731_ _1602_ _1604_ _1622_ _1624_ VPWR VGND sg13g2_or3_1
X_4662_ _1556_ mydesign.accum\[58\] _1558_ VPWR VGND sg13g2_xor2_1
XFILLER_31_1020 VPWR VGND sg13g2_decap_8
X_3613_ net626 VPWR _0635_ VGND mydesign.pe_inputs\[60\] net487 sg13g2_o21ai_1
X_4593_ _1483_ _1499_ _1480_ _1501_ VPWR VGND sg13g2_nand3_1
X_3544_ _0571_ _0557_ _0570_ VPWR VGND sg13g2_xnor2_1
X_3475_ VGND VPWR net554 mydesign.inputs\[0\]\[23\] _0510_ _0509_ sg13g2_a21oi_1
X_5214_ _2029_ _2045_ _2046_ VPWR VGND sg13g2_and2_1
X_5145_ _1968_ _1983_ _1965_ _1985_ VPWR VGND sg13g2_nand3_1
X_5076_ net475 VPWR _1920_ VGND net584 net913 sg13g2_o21ai_1
X_4027_ _1001_ _0999_ _1000_ VPWR VGND sg13g2_nand2_1
XFILLER_38_895 VPWR VGND sg13g2_decap_8
XFILLER_25_512 VPWR VGND sg13g2_fill_2
XFILLER_40_526 VPWR VGND sg13g2_decap_4
X_5978_ net201 VGND VPWR net691 mydesign.accum\[64\] clknet_leaf_40_clk sg13g2_dfrbpq_2
X_4929_ VGND VPWR net664 _1785_ _0260_ _1786_ sg13g2_a21oi_1
XFILLER_48_615 VPWR VGND sg13g2_decap_8
XFILLER_44_876 VPWR VGND sg13g2_decap_8
XFILLER_43_331 VPWR VGND sg13g2_decap_4
XFILLER_7_276 VPWR VGND sg13g2_fill_2
XFILLER_4_983 VPWR VGND sg13g2_decap_8
X_3260_ net775 _2670_ _2672_ _0028_ VPWR VGND sg13g2_mux2_1
X_3191_ net760 _2623_ net621 _2626_ VPWR VGND sg13g2_nand3_1
XFILLER_47_670 VPWR VGND sg13g2_decap_8
X_5901_ net351 VGND VPWR _0127_ mydesign.accum\[107\] clknet_leaf_41_clk sg13g2_dfrbpq_2
XFILLER_35_854 VPWR VGND sg13g2_fill_1
X_5832_ net105 VGND VPWR _0058_ mydesign.load_counter\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_2
XFILLER_35_887 VPWR VGND sg13g2_decap_8
X_5763_ net784 _2487_ _2510_ _0370_ VPWR VGND sg13g2_mux2_1
XFILLER_22_537 VPWR VGND sg13g2_decap_8
X_4714_ _1608_ _1585_ _1587_ VPWR VGND sg13g2_nand2_1
X_5694_ _2472_ _2473_ _0338_ VPWR VGND sg13g2_nor2_1
X_4645_ _1543_ net560 mydesign.pe_weights\[44\] _1521_ VPWR VGND sg13g2_and3_1
X_4576_ _1462_ VPWR _1485_ VGND _1461_ _1464_ sg13g2_o21ai_1
X_3527_ net467 VPWR _0555_ VGND net558 net958 sg13g2_o21ai_1
X_3458_ _0497_ net652 _0493_ VPWR VGND sg13g2_nand2_1
X_3389_ VGND VPWR _0405_ _0431_ _0437_ _2698_ sg13g2_a21oi_1
XFILLER_29_103 VPWR VGND sg13g2_fill_2
X_5128_ _1969_ _1964_ _1967_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_618 VPWR VGND sg13g2_decap_8
X_6017__398 VPWR VGND net398 sg13g2_tiehi
XFILLER_17_309 VPWR VGND sg13g2_decap_8
X_5059_ _1902_ _1901_ _1904_ VPWR VGND sg13g2_xor2_1
XFILLER_25_320 VPWR VGND sg13g2_fill_1
XFILLER_25_342 VPWR VGND sg13g2_decap_4
XFILLER_41_846 VPWR VGND sg13g2_decap_8
X_5807__139 VPWR VGND net139 sg13g2_tiehi
XFILLER_0_430 VPWR VGND sg13g2_decap_4
XFILLER_49_902 VPWR VGND sg13g2_decap_8
XFILLER_0_452 VPWR VGND sg13g2_decap_8
XFILLER_1_964 VPWR VGND sg13g2_decap_8
XFILLER_49_979 VPWR VGND sg13g2_decap_8
Xhold71 mydesign.accum\[64\] VPWR VGND net690 sg13g2_dlygate4sd3_1
Xhold82 mydesign.weights\[3\]\[6\] VPWR VGND net701 sg13g2_dlygate4sd3_1
Xhold60 mydesign.weights\[1\]\[17\] VPWR VGND net679 sg13g2_dlygate4sd3_1
Xhold93 mydesign.inputs\[3\]\[2\] VPWR VGND net712 sg13g2_dlygate4sd3_1
XFILLER_28_191 VPWR VGND sg13g2_decap_4
XFILLER_44_673 VPWR VGND sg13g2_decap_8
XFILLER_31_301 VPWR VGND sg13g2_fill_1
XFILLER_43_194 VPWR VGND sg13g2_decap_4
X_4430_ _1354_ _1355_ _1356_ VPWR VGND sg13g2_and2_1
X_6100_ net276 VGND VPWR net1041 mydesign.accum\[2\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_4361_ VGND VPWR _2558_ net441 _0185_ _1293_ sg13g2_a21oi_1
X_4292_ mydesign.pe_inputs\[45\] net539 mydesign.accum\[84\] _1234_ VPWR VGND sg13g2_a21o_1
X_3312_ _2696_ VPWR _0056_ VGND net597 net429 sg13g2_o21ai_1
Xfanout509 net510 net509 VPWR VGND sg13g2_buf_8
X_3243_ _2620_ net1109 _2663_ VPWR VGND sg13g2_nor2_1
X_6031_ net334 VGND VPWR net863 mydesign.pe_weights\[21\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3174_ _2611_ VPWR _0002_ VGND net432 _2612_ sg13g2_o21ai_1
X_6086__396 VPWR VGND net396 sg13g2_tiehi
XFILLER_22_334 VPWR VGND sg13g2_fill_2
X_5815_ net127 VGND VPWR _0041_ mydesign.inputs\[1\]\[20\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5746_ _2502_ VPWR _0361_ VGND _1771_ _2500_ sg13g2_o21ai_1
X_5677_ _2462_ VPWR _0332_ VGND net604 _2461_ sg13g2_o21ai_1
X_4628_ net625 VPWR _1532_ VGND net1090 net438 sg13g2_o21ai_1
X_4559_ _1468_ VPWR _1469_ VGND _1447_ _1449_ sg13g2_o21ai_1
XFILLER_14_802 VPWR VGND sg13g2_fill_2
XFILLER_41_643 VPWR VGND sg13g2_fill_1
XFILLER_41_698 VPWR VGND sg13g2_fill_1
XFILLER_1_794 VPWR VGND sg13g2_decap_8
XFILLER_49_776 VPWR VGND sg13g2_decap_8
XFILLER_37_938 VPWR VGND sg13g2_decap_8
X_6070__186 VPWR VGND net186 sg13g2_tiehi
XFILLER_45_982 VPWR VGND sg13g2_decap_8
X_3930_ net459 VPWR _0912_ VGND mydesign.weights\[3\]\[8\] net547 sg13g2_o21ai_1
XFILLER_16_150 VPWR VGND sg13g2_fill_1
X_3861_ _0852_ _0835_ _0850_ VPWR VGND sg13g2_xnor2_1
X_5600_ _2391_ mydesign.pe_inputs\[6\] mydesign.pe_weights\[17\] VPWR VGND sg13g2_nand2_1
X_3792_ _0788_ VPWR _0789_ VGND _0785_ _0786_ sg13g2_o21ai_1
X_5531_ _2331_ VPWR _2332_ VGND net592 net1089 sg13g2_o21ai_1
XFILLER_8_360 VPWR VGND sg13g2_decap_4
X_5462_ _2264_ _2261_ _2266_ VPWR VGND sg13g2_xor2_1
X_5393_ net481 VPWR _2207_ VGND net590 net1042 sg13g2_o21ai_1
X_4413_ _1340_ _1324_ _1338_ VPWR VGND sg13g2_xnor2_1
X_4344_ _1268_ VPWR _1283_ VGND _1267_ _1271_ sg13g2_o21ai_1
X_4275_ _1196_ _1217_ _1218_ VPWR VGND sg13g2_nor2b_1
X_6014_ net34 VGND VPWR _0240_ mydesign.accum\[52\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3226_ net623 _2649_ _2650_ VPWR VGND sg13g2_and2_1
X_3157_ net756 net744 _2584_ _2598_ VPWR VGND sg13g2_nand3_1
X_5914__329 VPWR VGND net329 sg13g2_tiehi
XFILLER_27_404 VPWR VGND sg13g2_decap_8
XFILLER_28_949 VPWR VGND sg13g2_decap_8
X_3088_ VPWR _2529_ net816 VGND sg13g2_inv_1
XFILLER_36_993 VPWR VGND sg13g2_decap_8
XFILLER_10_326 VPWR VGND sg13g2_decap_8
X_5729_ net711 _2490_ net615 _2493_ VPWR VGND sg13g2_nand3_1
Xhold360 mydesign.accum\[24\] VPWR VGND net979 sg13g2_dlygate4sd3_1
Xhold371 mydesign.accum\[59\] VPWR VGND net990 sg13g2_dlygate4sd3_1
Xhold393 mydesign.accum\[28\] VPWR VGND net1012 sg13g2_dlygate4sd3_1
Xhold382 _0299_ VPWR VGND net1001 sg13g2_dlygate4sd3_1
XFILLER_19_927 VPWR VGND sg13g2_decap_8
XFILLER_46_768 VPWR VGND sg13g2_decap_8
XFILLER_26_470 VPWR VGND sg13g2_decap_8
X_5965__227 VPWR VGND net227 sg13g2_tiehi
XFILLER_42_996 VPWR VGND sg13g2_decap_8
XFILLER_41_484 VPWR VGND sg13g2_fill_2
XFILLER_14_698 VPWR VGND sg13g2_fill_1
XFILLER_3_32 VPWR VGND sg13g2_fill_1
XFILLER_49_540 VPWR VGND sg13g2_decap_8
X_4060_ _1016_ _1031_ _1008_ _1032_ VPWR VGND sg13g2_nand3_1
XFILLER_3_1027 VPWR VGND sg13g2_fill_2
XFILLER_18_960 VPWR VGND sg13g2_decap_8
XFILLER_24_418 VPWR VGND sg13g2_decap_8
X_4962_ net531 net528 mydesign.accum\[43\] _1817_ VPWR VGND sg13g2_nand3_1
X_4893_ _1765_ net671 _1762_ VPWR VGND sg13g2_nand2_1
X_3913_ _0901_ _0885_ _0899_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_952 VPWR VGND sg13g2_decap_8
X_3844_ _0827_ VPWR _0835_ VGND _0808_ _0825_ sg13g2_o21ai_1
XFILLER_20_646 VPWR VGND sg13g2_decap_4
X_3775_ net628 VPWR _0776_ VGND net1024 net433 sg13g2_o21ai_1
XFILLER_9_691 VPWR VGND sg13g2_fill_2
X_5514_ VGND VPWR net592 _2314_ _0316_ _2315_ sg13g2_a21oi_1
X_5445_ _2250_ mydesign.accum\[9\] net521 mydesign.pe_weights\[21\] VPWR VGND sg13g2_and3_2
X_5376_ _2190_ mydesign.pe_inputs\[14\] mydesign.pe_weights\[26\] VPWR VGND sg13g2_nand2_1
X_4327_ VGND VPWR net539 mydesign.pe_inputs\[47\] _1267_ mydesign.accum\[86\] sg13g2_a21oi_1
X_4258_ _1184_ _1200_ _1202_ VPWR VGND sg13g2_nor2_1
XFILLER_41_1000 VPWR VGND sg13g2_decap_8
X_3209_ _2637_ VPWR _0012_ VGND _2517_ _2633_ sg13g2_o21ai_1
X_6131__356 VPWR VGND net356 sg13g2_tiehi
X_4189_ VGND VPWR mydesign.accum\[92\] _1124_ _1146_ _1126_ sg13g2_a21oi_1
XFILLER_43_705 VPWR VGND sg13g2_fill_2
XFILLER_24_930 VPWR VGND sg13g2_decap_8
XFILLER_24_974 VPWR VGND sg13g2_decap_8
XFILLER_3_823 VPWR VGND sg13g2_decap_8
XFILLER_2_311 VPWR VGND sg13g2_decap_8
XFILLER_2_322 VPWR VGND sg13g2_fill_2
XFILLER_3_889 VPWR VGND sg13g2_fill_2
Xhold190 _0084_ VPWR VGND net809 sg13g2_dlygate4sd3_1
XFILLER_27_790 VPWR VGND sg13g2_decap_8
XFILLER_33_204 VPWR VGND sg13g2_decap_8
XFILLER_33_215 VPWR VGND sg13g2_fill_1
XFILLER_18_1002 VPWR VGND sg13g2_decap_8
XFILLER_30_955 VPWR VGND sg13g2_decap_8
X_5785__167 VPWR VGND net167 sg13g2_tiehi
X_3560_ _0586_ _0580_ _0585_ VPWR VGND sg13g2_nand2_1
XFILLER_5_182 VPWR VGND sg13g2_decap_8
X_5230_ _2059_ _2060_ _2036_ _2061_ VPWR VGND sg13g2_nand3_1
X_3491_ _2586_ _0522_ _0523_ VPWR VGND sg13g2_and2_1
X_5161_ mydesign.inputs\[3\]\[4\] net549 _1999_ VPWR VGND sg13g2_nor2b_1
X_4112_ _1073_ net808 _1051_ VPWR VGND sg13g2_nand2_1
X_5092_ _1935_ _1911_ _1933_ VPWR VGND sg13g2_xnor2_1
X_4043_ _1014_ _1013_ _1016_ VPWR VGND sg13g2_xor2_1
XFILLER_49_370 VPWR VGND sg13g2_decap_4
X_5994_ net134 VGND VPWR net687 mydesign.accum\[56\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_4945_ _1801_ _1799_ _1800_ VPWR VGND sg13g2_nand2_1
X_4876_ _1750_ VPWR _1752_ VGND _1737_ _1740_ sg13g2_o21ai_1
X_3827_ VGND VPWR _0793_ _0795_ _0819_ _2583_ sg13g2_a21oi_1
XFILLER_21_988 VPWR VGND sg13g2_decap_8
X_3758_ _0764_ net973 _0765_ VPWR VGND sg13g2_xor2_1
XFILLER_20_498 VPWR VGND sg13g2_fill_2
X_3689_ _0698_ _0699_ _0678_ _0700_ VPWR VGND sg13g2_nand3_1
X_5428_ VGND VPWR _2215_ _2230_ _2239_ _2229_ sg13g2_a21oi_1
X_5359_ _2174_ _2172_ _2173_ VPWR VGND sg13g2_nand2_1
XFILLER_0_859 VPWR VGND sg13g2_decap_8
XFILLER_28_532 VPWR VGND sg13g2_decap_4
XFILLER_43_524 VPWR VGND sg13g2_decap_4
XFILLER_24_793 VPWR VGND sg13g2_fill_2
XFILLER_12_977 VPWR VGND sg13g2_decap_8
XFILLER_11_487 VPWR VGND sg13g2_fill_1
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_697 VPWR VGND sg13g2_fill_1
XFILLER_17_7 VPWR VGND sg13g2_fill_1
XFILLER_47_852 VPWR VGND sg13g2_decap_8
XFILLER_34_557 VPWR VGND sg13g2_fill_2
X_4730_ _1622_ VPWR _1623_ VGND _1602_ _1604_ sg13g2_o21ai_1
XFILLER_9_86 VPWR VGND sg13g2_fill_1
XFILLER_30_774 VPWR VGND sg13g2_fill_2
X_4661_ mydesign.pe_weights\[46\] _1521_ mydesign.accum\[58\] _1557_ VPWR VGND sg13g2_nand3_1
X_3612_ VGND VPWR net559 _0633_ _0095_ _0634_ sg13g2_a21oi_1
X_4592_ VGND VPWR _1480_ _1483_ _1500_ _1499_ sg13g2_a21oi_1
X_3543_ _0567_ _0545_ _0570_ VPWR VGND sg13g2_xor2_1
XFILLER_7_981 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
X_3474_ net554 mydesign.inputs\[0\]\[27\] _0509_ VPWR VGND sg13g2_nor2b_1
X_5213_ _2045_ _2035_ _2043_ VPWR VGND sg13g2_xnor2_1
X_5144_ VGND VPWR _1965_ _1968_ _1984_ _1983_ sg13g2_a21oi_1
X_5878__393 VPWR VGND net393 sg13g2_tiehi
XFILLER_38_841 VPWR VGND sg13g2_decap_4
X_5075_ _1919_ _1903_ _1918_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_329 VPWR VGND sg13g2_decap_8
XFILLER_38_874 VPWR VGND sg13g2_decap_8
X_4026_ _0977_ _0953_ _0980_ _1000_ VPWR VGND sg13g2_a21o_1
XFILLER_44_17 VPWR VGND sg13g2_decap_8
XFILLER_25_557 VPWR VGND sg13g2_fill_1
X_5977_ net203 VGND VPWR _0203_ mydesign.pe_weights\[35\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_4928_ net477 VPWR _1786_ VGND net664 _1785_ sg13g2_o21ai_1
X_4859_ _1736_ _1725_ _1734_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
X_6120__76 VPWR VGND net76 sg13g2_tiehi
XFILLER_18_62 VPWR VGND sg13g2_fill_2
XFILLER_43_310 VPWR VGND sg13g2_fill_1
XFILLER_18_95 VPWR VGND sg13g2_decap_8
XFILLER_29_885 VPWR VGND sg13g2_decap_8
XFILLER_44_855 VPWR VGND sg13g2_decap_8
XFILLER_7_222 VPWR VGND sg13g2_fill_2
XFILLER_12_796 VPWR VGND sg13g2_fill_2
XFILLER_4_962 VPWR VGND sg13g2_decap_8
X_3190_ _2624_ VPWR _0005_ VGND _2623_ net603 sg13g2_o21ai_1
XFILLER_39_649 VPWR VGND sg13g2_fill_2
X_5900_ net353 VGND VPWR net1011 mydesign.accum\[106\] clknet_leaf_41_clk sg13g2_dfrbpq_2
X_5831_ net107 VGND VPWR _0057_ mydesign.load_counter\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_2
X_5762_ net803 _2486_ _2510_ _0369_ VPWR VGND sg13g2_mux2_1
X_4713_ _1605_ _1594_ _1607_ VPWR VGND sg13g2_xor2_1
X_5693_ VGND VPWR net457 _2467_ _2473_ net512 sg13g2_a21oi_1
X_4644_ VGND VPWR _2549_ net437 _0219_ _1542_ sg13g2_a21oi_1
XFILLER_30_593 VPWR VGND sg13g2_fill_1
X_4575_ _1482_ _1479_ _1484_ VPWR VGND sg13g2_xor2_1
X_3526_ _0554_ _0537_ _0552_ VPWR VGND sg13g2_xnor2_1
X_3457_ _0496_ VPWR _0078_ VGND net599 _0492_ sg13g2_o21ai_1
X_3388_ VGND VPWR net504 _0434_ _0436_ _0435_ sg13g2_a21oi_1
X_5127_ VGND VPWR _1968_ _1967_ _1964_ sg13g2_or2_1
X_5058_ mydesign.pe_weights\[32\] net1107 net734 _1903_ VPWR VGND _1901_ sg13g2_nand4_1
X_4009_ _0982_ _0983_ _0984_ VPWR VGND sg13g2_nor2b_1
X_5924__309 VPWR VGND net309 sg13g2_tiehi
XFILLER_4_236 VPWR VGND sg13g2_fill_1
XFILLER_20_85 VPWR VGND sg13g2_decap_8
XFILLER_1_943 VPWR VGND sg13g2_decap_8
X_5900__353 VPWR VGND net353 sg13g2_tiehi
XFILLER_49_958 VPWR VGND sg13g2_decap_8
XFILLER_48_435 VPWR VGND sg13g2_fill_2
XFILLER_0_486 VPWR VGND sg13g2_fill_2
Xhold50 mydesign.inputs\[2\]\[7\] VPWR VGND net669 sg13g2_dlygate4sd3_1
XFILLER_48_468 VPWR VGND sg13g2_fill_1
Xhold72 _0204_ VPWR VGND net691 sg13g2_dlygate4sd3_1
Xhold83 _0114_ VPWR VGND net702 sg13g2_dlygate4sd3_1
Xhold61 mydesign.inputs\[3\]\[11\] VPWR VGND net680 sg13g2_dlygate4sd3_1
Xhold94 _0055_ VPWR VGND net713 sg13g2_dlygate4sd3_1
XFILLER_29_660 VPWR VGND sg13g2_fill_2
XFILLER_17_866 VPWR VGND sg13g2_fill_1
XFILLER_44_652 VPWR VGND sg13g2_decap_8
XFILLER_16_343 VPWR VGND sg13g2_fill_1
XFILLER_32_869 VPWR VGND sg13g2_fill_1
XFILLER_8_520 VPWR VGND sg13g2_decap_8
XFILLER_31_379 VPWR VGND sg13g2_decap_8
X_4360_ net633 VPWR _1293_ VGND net862 net441 sg13g2_o21ai_1
X_5975__207 VPWR VGND net207 sg13g2_tiehi
X_3311_ net719 net429 net618 _2696_ VPWR VGND sg13g2_nand3_1
X_4291_ net539 mydesign.pe_inputs\[45\] mydesign.accum\[84\] _1233_ VPWR VGND sg13g2_nand3_1
XFILLER_3_280 VPWR VGND sg13g2_fill_1
X_6030_ net342 VGND VPWR _0256_ mydesign.pe_weights\[20\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3242_ _2662_ net614 net605 VPWR VGND sg13g2_nand2_1
XFILLER_6_1014 VPWR VGND sg13g2_decap_8
X_3173_ _2612_ net733 net616 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_46_clk clknet_3_1__leaf_clk clknet_leaf_46_clk VPWR VGND sg13g2_buf_8
XFILLER_35_674 VPWR VGND sg13g2_fill_1
X_5814_ net128 VGND VPWR _0040_ mydesign.inputs\[1\]\[19\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_35_696 VPWR VGND sg13g2_decap_4
XFILLER_10_508 VPWR VGND sg13g2_decap_4
X_5745_ _2502_ net727 _2500_ VPWR VGND sg13g2_nand2_1
XFILLER_30_390 VPWR VGND sg13g2_fill_1
X_5676_ _2462_ net683 _2461_ VPWR VGND sg13g2_nand2_1
X_6023__370 VPWR VGND net370 sg13g2_tiehi
X_4627_ _1531_ _1530_ _0392_ _1529_ net460 VPWR VGND sg13g2_a22oi_1
X_4558_ _1467_ _1459_ _1468_ VPWR VGND sg13g2_xor2_1
X_4489_ net633 VPWR _1407_ VGND mydesign.pe_weights\[48\] net491 sg13g2_o21ai_1
X_3509_ _0536_ _0535_ _0538_ VPWR VGND sg13g2_xor2_1
XFILLER_18_608 VPWR VGND sg13g2_decap_8
XFILLER_39_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_37_clk clknet_3_5__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_41_666 VPWR VGND sg13g2_fill_2
XFILLER_5_523 VPWR VGND sg13g2_fill_2
XFILLER_5_512 VPWR VGND sg13g2_decap_8
XFILLER_12_1019 VPWR VGND sg13g2_decap_8
XFILLER_5_545 VPWR VGND sg13g2_fill_2
XFILLER_49_755 VPWR VGND sg13g2_decap_8
XFILLER_37_917 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_28_clk clknet_3_7__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_45_961 VPWR VGND sg13g2_decap_8
XFILLER_17_652 VPWR VGND sg13g2_fill_1
X_5840__89 VPWR VGND net89 sg13g2_tiehi
X_3860_ _0851_ _0835_ _0850_ VPWR VGND sg13g2_nand2_1
X_3791_ _0788_ _0392_ _0787_ VPWR VGND sg13g2_nand2_1
XFILLER_32_699 VPWR VGND sg13g2_decap_4
X_5530_ net592 VPWR _2331_ VGND _2329_ _2330_ sg13g2_o21ai_1
X_5461_ _2261_ _2264_ _2265_ VPWR VGND sg13g2_nor2_1
X_6002__86 VPWR VGND net86 sg13g2_tiehi
X_4412_ _1324_ _1338_ _1339_ VPWR VGND sg13g2_and2_1
X_5392_ VGND VPWR _2204_ _2205_ _2206_ net503 sg13g2_a21oi_1
X_4343_ _1282_ _1276_ _1279_ VPWR VGND sg13g2_nand2_1
XFILLER_28_1026 VPWR VGND sg13g2_fill_2
X_4274_ _1216_ _1213_ _1217_ VPWR VGND sg13g2_xor2_1
X_3225_ _2638_ _2647_ net605 _2649_ VPWR VGND sg13g2_nand3_1
X_6013_ net38 VGND VPWR _0239_ mydesign.accum\[51\] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_39_221 VPWR VGND sg13g2_fill_1
X_3156_ _2597_ net541 net496 VPWR VGND sg13g2_nand2_1
XFILLER_28_928 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_19_clk clknet_3_3__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
X_3087_ VPWR _2528_ net773 VGND sg13g2_inv_1
XFILLER_36_972 VPWR VGND sg13g2_decap_8
XFILLER_35_460 VPWR VGND sg13g2_fill_2
X_3989_ VGND VPWR _0939_ _0955_ _0964_ _0957_ sg13g2_a21oi_1
X_5728_ _2492_ VPWR _0353_ VGND net602 _2490_ sg13g2_o21ai_1
X_5659_ _2447_ net519 mydesign.pe_weights\[19\] _2446_ VPWR VGND sg13g2_and3_1
XFILLER_7_6 VPWR VGND sg13g2_fill_1
Xhold361 mydesign.accum\[47\] VPWR VGND net980 sg13g2_dlygate4sd3_1
Xhold350 mydesign.accum\[51\] VPWR VGND net969 sg13g2_dlygate4sd3_1
Xhold383 mydesign.accum\[36\] VPWR VGND net1002 sg13g2_dlygate4sd3_1
Xhold394 mydesign.pe_weights\[40\] VPWR VGND net1013 sg13g2_dlygate4sd3_1
Xhold372 mydesign.accum\[112\] VPWR VGND net991 sg13g2_dlygate4sd3_1
XFILLER_46_747 VPWR VGND sg13g2_decap_8
XFILLER_27_983 VPWR VGND sg13g2_decap_8
XFILLER_42_975 VPWR VGND sg13g2_decap_8
XFILLER_41_441 VPWR VGND sg13g2_decap_8
XFILLER_41_430 VPWR VGND sg13g2_fill_1
XFILLER_13_121 VPWR VGND sg13g2_fill_2
XFILLER_26_95 VPWR VGND sg13g2_decap_4
XFILLER_10_861 VPWR VGND sg13g2_decap_4
XFILLER_6_876 VPWR VGND sg13g2_fill_1
XFILLER_47_7 VPWR VGND sg13g2_fill_2
XFILLER_3_1006 VPWR VGND sg13g2_decap_8
XFILLER_24_408 VPWR VGND sg13g2_fill_1
XFILLER_17_460 VPWR VGND sg13g2_fill_1
X_4961_ _1816_ mydesign.pe_weights\[38\] mydesign.pe_inputs\[25\] VPWR VGND sg13g2_nand2_1
XFILLER_33_931 VPWR VGND sg13g2_decap_8
XFILLER_44_290 VPWR VGND sg13g2_decap_4
X_4892_ _1764_ VPWR _0245_ VGND net601 _1761_ sg13g2_o21ai_1
X_3912_ _0885_ _0899_ _0900_ VPWR VGND sg13g2_nor2b_1
X_3843_ _0829_ _0831_ _0834_ VPWR VGND sg13g2_and2_1
X_3774_ VGND VPWR _2583_ net433 _0116_ _0775_ sg13g2_a21oi_1
X_5513_ net481 VPWR _2315_ VGND net592 net1048 sg13g2_o21ai_1
X_5444_ VGND VPWR net729 _2248_ _0312_ _2249_ sg13g2_a21oi_1
Xclkbuf_leaf_8_clk clknet_3_3__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_5375_ _2172_ VPWR _2189_ VGND _2171_ _2174_ sg13g2_o21ai_1
X_4326_ _1266_ _1265_ _0177_ VPWR VGND sg13g2_nor2b_1
X_4257_ _1201_ _1184_ _1200_ VPWR VGND sg13g2_nand2_1
X_4188_ _1145_ _1141_ _1143_ VPWR VGND sg13g2_xnor2_1
X_3208_ net617 _2633_ net662 _2637_ VPWR VGND sg13g2_nand3_1
X_3139_ VPWR _2580_ net1046 VGND sg13g2_inv_1
XFILLER_27_224 VPWR VGND sg13g2_fill_1
XFILLER_27_246 VPWR VGND sg13g2_decap_8
XFILLER_43_739 VPWR VGND sg13g2_decap_8
XFILLER_24_953 VPWR VGND sg13g2_decap_8
XFILLER_23_452 VPWR VGND sg13g2_fill_1
XFILLER_10_135 VPWR VGND sg13g2_fill_2
XFILLER_10_168 VPWR VGND sg13g2_fill_2
XFILLER_12_75 VPWR VGND sg13g2_fill_1
Xhold180 mydesign.inputs\[1\]\[9\] VPWR VGND net799 sg13g2_dlygate4sd3_1
Xhold191 mydesign.weights\[2\]\[14\] VPWR VGND net810 sg13g2_dlygate4sd3_1
XFILLER_18_257 VPWR VGND sg13g2_fill_2
XFILLER_34_728 VPWR VGND sg13g2_fill_2
XFILLER_14_474 VPWR VGND sg13g2_fill_2
XFILLER_15_986 VPWR VGND sg13g2_decap_8
XFILLER_41_282 VPWR VGND sg13g2_fill_2
XFILLER_14_485 VPWR VGND sg13g2_fill_2
XFILLER_30_934 VPWR VGND sg13g2_decap_8
X_3490_ net553 mydesign.weights\[0\]\[26\] mydesign.weights\[0\]\[22\] mydesign.weights\[0\]\[18\]
+ mydesign.weights\[0\]\[14\] net546 _0522_ VPWR VGND sg13g2_mux4_1
XFILLER_6_673 VPWR VGND sg13g2_fill_1
X_5160_ VGND VPWR net575 _1997_ _0279_ _1998_ sg13g2_a21oi_1
X_4111_ _1072_ _1070_ _1071_ VPWR VGND sg13g2_nand2_1
X_5091_ _1934_ _1911_ _1933_ VPWR VGND sg13g2_nand2_1
X_4042_ _1015_ _1013_ _1014_ VPWR VGND sg13g2_nand2_1
XFILLER_37_522 VPWR VGND sg13g2_fill_2
XFILLER_37_511 VPWR VGND sg13g2_decap_8
X_5833__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_37_599 VPWR VGND sg13g2_decap_8
X_5993_ net138 VGND VPWR _0219_ mydesign.pe_weights\[31\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_4944_ net528 mydesign.pe_weights\[38\] mydesign.accum\[42\] _1800_ VPWR VGND sg13g2_a21o_1
X_4875_ _1737_ _1740_ _1750_ _1751_ VPWR VGND sg13g2_or3_1
X_3826_ _0818_ mydesign.pe_inputs\[58\] _0783_ VPWR VGND sg13g2_nand2_1
XFILLER_21_967 VPWR VGND sg13g2_decap_8
X_3757_ _0748_ VPWR _0764_ VGND _0747_ _0751_ sg13g2_o21ai_1
X_3688_ _0690_ VPWR _0699_ VGND _0696_ _0697_ sg13g2_o21ai_1
X_5868__37 VPWR VGND net37 sg13g2_tiehi
X_5427_ _2235_ VPWR _2238_ VGND _2218_ _2231_ sg13g2_o21ai_1
XFILLER_0_838 VPWR VGND sg13g2_decap_8
X_5358_ net527 mydesign.pe_inputs\[12\] mydesign.accum\[19\] _2173_ VPWR VGND sg13g2_a21o_1
X_4309_ _1250_ mydesign.pe_weights\[58\] mydesign.pe_inputs\[47\] VPWR VGND sg13g2_nand2_1
XFILLER_47_308 VPWR VGND sg13g2_fill_2
X_5289_ _2117_ _2116_ _2102_ VPWR VGND sg13g2_nand2b_1
XFILLER_12_912 VPWR VGND sg13g2_decap_4
XFILLER_12_956 VPWR VGND sg13g2_decap_8
XFILLER_48_1007 VPWR VGND sg13g2_decap_8
XFILLER_3_610 VPWR VGND sg13g2_fill_1
XFILLER_3_654 VPWR VGND sg13g2_fill_2
XFILLER_3_0 VPWR VGND sg13g2_fill_1
XFILLER_3_676 VPWR VGND sg13g2_fill_2
XFILLER_47_831 VPWR VGND sg13g2_decap_8
Xfanout490 _2602_ net490 VPWR VGND sg13g2_buf_8
XFILLER_46_352 VPWR VGND sg13g2_fill_1
XFILLER_34_514 VPWR VGND sg13g2_decap_4
X_4660_ mydesign.pe_weights\[46\] VPWR _1556_ VGND _1517_ _1520_ sg13g2_o21ai_1
X_3611_ net468 VPWR _0634_ VGND net559 net1004 sg13g2_o21ai_1
X_4591_ _1499_ _1497_ _1498_ VPWR VGND sg13g2_nand2_1
X_3542_ _0545_ _0567_ _0569_ VPWR VGND sg13g2_nor2_1
X_3473_ _0507_ _0508_ _0082_ VPWR VGND sg13g2_nor2_1
XFILLER_6_492 VPWR VGND sg13g2_fill_2
XFILLER_9_1012 VPWR VGND sg13g2_decap_8
X_5212_ _2044_ _2043_ _2035_ VPWR VGND sg13g2_nand2b_1
X_5143_ _1983_ _1981_ _1982_ VPWR VGND sg13g2_nand2_1
XFILLER_36_0 VPWR VGND sg13g2_decap_4
XFILLER_29_308 VPWR VGND sg13g2_decap_8
X_5074_ _1918_ _1899_ _1916_ VPWR VGND sg13g2_xnor2_1
X_4025_ _0999_ _0987_ _0997_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_330 VPWR VGND sg13g2_decap_4
XFILLER_25_514 VPWR VGND sg13g2_fill_1
X_5976_ net205 VGND VPWR _0202_ mydesign.pe_weights\[34\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_4927_ net501 _2536_ _2540_ _1785_ VPWR VGND sg13g2_nor3_1
X_4858_ _1735_ _1725_ _1734_ VPWR VGND sg13g2_nand2_1
XFILLER_21_742 VPWR VGND sg13g2_fill_2
XFILLER_21_753 VPWR VGND sg13g2_fill_2
X_3809_ VGND VPWR _0804_ _0803_ _0800_ sg13g2_or2_1
XFILLER_20_263 VPWR VGND sg13g2_decap_4
XFILLER_5_908 VPWR VGND sg13g2_decap_8
X_4789_ _1669_ mydesign.pe_weights\[41\] mydesign.pe_inputs\[29\] VPWR VGND sg13g2_nand2_1
XFILLER_4_429 VPWR VGND sg13g2_fill_1
XFILLER_4_418 VPWR VGND sg13g2_decap_8
XFILLER_0_613 VPWR VGND sg13g2_decap_8
XFILLER_0_657 VPWR VGND sg13g2_decap_8
X_5892__369 VPWR VGND net369 sg13g2_tiehi
XFILLER_29_831 VPWR VGND sg13g2_decap_4
XFILLER_44_834 VPWR VGND sg13g2_decap_8
XFILLER_29_875 VPWR VGND sg13g2_fill_1
XFILLER_43_344 VPWR VGND sg13g2_fill_2
XFILLER_28_396 VPWR VGND sg13g2_fill_1
XFILLER_43_377 VPWR VGND sg13g2_decap_8
XFILLER_15_1028 VPWR VGND sg13g2_fill_1
Xheichips25_template_400 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_11_263 VPWR VGND sg13g2_fill_2
XFILLER_7_278 VPWR VGND sg13g2_fill_1
XFILLER_3_462 VPWR VGND sg13g2_decap_8
XFILLER_3_440 VPWR VGND sg13g2_decap_4
XFILLER_3_473 VPWR VGND sg13g2_fill_2
X_6149__256 VPWR VGND net256 sg13g2_tiehi
X_5830_ net109 VGND VPWR net720 mydesign.inputs\[3\]\[3\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_5761_ net767 _2485_ _2510_ _0368_ VPWR VGND sg13g2_mux2_1
XFILLER_30_550 VPWR VGND sg13g2_fill_1
X_4712_ _1606_ _1605_ _1594_ VPWR VGND sg13g2_nand2b_1
X_5692_ _2466_ _2471_ _2472_ VPWR VGND sg13g2_nor2_1
X_4643_ net625 VPWR _1542_ VGND net1077 net437 sg13g2_o21ai_1
X_4574_ VGND VPWR _1483_ _1482_ _1479_ sg13g2_or2_1
X_3525_ VGND VPWR _0553_ _0552_ _0537_ sg13g2_or2_1
X_3456_ _0496_ net418 _0493_ VPWR VGND sg13g2_nand2_1
X_3387_ net457 VPWR _0435_ VGND net504 _0432_ sg13g2_o21ai_1
X_5126_ _1967_ _1965_ _1966_ VPWR VGND sg13g2_nand2_1
XFILLER_45_609 VPWR VGND sg13g2_fill_1
X_5057_ mydesign.pe_weights\[32\] net526 net734 _1902_ VPWR VGND sg13g2_nand3_1
X_4008_ _0964_ VPWR _0983_ VGND _0980_ _0981_ sg13g2_o21ai_1
XFILLER_38_694 VPWR VGND sg13g2_fill_1
XFILLER_25_311 VPWR VGND sg13g2_decap_8
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
XFILLER_13_528 VPWR VGND sg13g2_fill_1
X_5959_ net239 VGND VPWR _0185_ mydesign.pe_weights\[37\] clknet_leaf_41_clk sg13g2_dfrbpq_2
XFILLER_21_583 VPWR VGND sg13g2_fill_2
XFILLER_21_594 VPWR VGND sg13g2_decap_8
XFILLER_20_31 VPWR VGND sg13g2_fill_2
XFILLER_1_922 VPWR VGND sg13g2_decap_8
XFILLER_49_937 VPWR VGND sg13g2_decap_8
XFILLER_0_465 VPWR VGND sg13g2_decap_8
XFILLER_1_999 VPWR VGND sg13g2_decap_8
Xhold40 _0321_ VPWR VGND net659 sg13g2_dlygate4sd3_1
X_5837__95 VPWR VGND net95 sg13g2_tiehi
Xhold62 _0323_ VPWR VGND net681 sg13g2_dlygate4sd3_1
Xhold73 mydesign.weights\[2\]\[18\] VPWR VGND net692 sg13g2_dlygate4sd3_1
Xhold51 mydesign.inputs\[2\]\[16\] VPWR VGND net670 sg13g2_dlygate4sd3_1
Xhold84 mydesign.inputs\[2\]\[18\] VPWR VGND net703 sg13g2_dlygate4sd3_1
Xhold95 mydesign.weights\[0\]\[27\] VPWR VGND net714 sg13g2_dlygate4sd3_1
XFILLER_29_650 VPWR VGND sg13g2_fill_1
XFILLER_44_631 VPWR VGND sg13g2_decap_8
XFILLER_17_834 VPWR VGND sg13g2_fill_1
XFILLER_43_174 VPWR VGND sg13g2_fill_1
XFILLER_12_561 VPWR VGND sg13g2_fill_1
XFILLER_8_554 VPWR VGND sg13g2_decap_8
XFILLER_4_771 VPWR VGND sg13g2_decap_4
X_3310_ _2695_ VPWR _0055_ VGND net599 net429 sg13g2_o21ai_1
X_4290_ _1232_ mydesign.pe_weights\[58\] mydesign.pe_inputs\[46\] VPWR VGND sg13g2_nand2_1
X_3241_ _2661_ net617 _2591_ VPWR VGND sg13g2_nand2_2
XFILLER_39_414 VPWR VGND sg13g2_fill_2
XFILLER_39_403 VPWR VGND sg13g2_decap_8
X_3172_ _2611_ net2 net432 VPWR VGND sg13g2_nand2_1
XFILLER_39_469 VPWR VGND sg13g2_decap_4
XFILLER_39_458 VPWR VGND sg13g2_fill_2
XFILLER_47_491 VPWR VGND sg13g2_fill_2
XFILLER_19_182 VPWR VGND sg13g2_fill_2
X_5813_ net129 VGND VPWR _0039_ mydesign.inputs\[1\]\[18\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_22_303 VPWR VGND sg13g2_fill_2
XFILLER_34_185 VPWR VGND sg13g2_fill_1
XFILLER_22_336 VPWR VGND sg13g2_fill_1
XFILLER_41_19 VPWR VGND sg13g2_decap_8
X_5744_ _2501_ VPWR _0360_ VGND _1769_ _2500_ sg13g2_o21ai_1
X_5675_ _2461_ net462 _2684_ VPWR VGND sg13g2_nand2_2
X_4626_ mydesign.inputs\[2\]\[18\] mydesign.inputs\[2\]\[14\] net557 _1530_ VPWR VGND
+ sg13g2_mux2_1
X_5806__141 VPWR VGND net141 sg13g2_tiehi
X_4557_ _1467_ _1460_ _1465_ VPWR VGND sg13g2_xnor2_1
X_4488_ _1406_ VPWR _0199_ VGND net597 _1401_ sg13g2_o21ai_1
X_3508_ net455 _0517_ net721 _0537_ VPWR VGND _0535_ sg13g2_nand4_1
X_3439_ net513 mydesign.accum\[103\] mydesign.accum\[71\] mydesign.accum\[39\] mydesign.accum\[7\]
+ net506 _0482_ VPWR VGND sg13g2_mux4_1
X_5109_ _1951_ _1943_ _1949_ VPWR VGND sg13g2_xnor2_1
Xheichips25_template_20 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_46_929 VPWR VGND sg13g2_decap_8
XFILLER_39_970 VPWR VGND sg13g2_decap_8
X_6089_ net368 VGND VPWR _0315_ mydesign.accum\[11\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_38_491 VPWR VGND sg13g2_fill_1
X_6030__342 VPWR VGND net342 sg13g2_tiehi
XFILLER_14_804 VPWR VGND sg13g2_fill_1
XFILLER_41_623 VPWR VGND sg13g2_decap_8
XFILLER_40_122 VPWR VGND sg13g2_decap_8
XFILLER_14_859 VPWR VGND sg13g2_fill_2
XFILLER_41_678 VPWR VGND sg13g2_decap_4
XFILLER_40_166 VPWR VGND sg13g2_decap_4
XFILLER_5_557 VPWR VGND sg13g2_decap_4
XFILLER_49_734 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_fill_2
XFILLER_45_940 VPWR VGND sg13g2_decap_8
XFILLER_16_141 VPWR VGND sg13g2_fill_1
XFILLER_17_686 VPWR VGND sg13g2_decap_8
XFILLER_32_623 VPWR VGND sg13g2_decap_8
XFILLER_32_634 VPWR VGND sg13g2_fill_2
X_3790_ mydesign.weights\[2\]\[17\] mydesign.weights\[2\]\[13\] net551 _0787_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_20_818 VPWR VGND sg13g2_decap_4
X_5460_ _2264_ _2262_ _2263_ VPWR VGND sg13g2_nand2_1
X_4411_ _1337_ _1325_ _1338_ VPWR VGND sg13g2_xor2_1
X_5391_ _2203_ VPWR _2205_ VGND _2183_ _2185_ sg13g2_o21ai_1
X_4342_ VGND VPWR net579 _1280_ _0178_ _1281_ sg13g2_a21oi_1
XFILLER_28_1005 VPWR VGND sg13g2_decap_8
X_4273_ _1216_ _1214_ _1215_ VPWR VGND sg13g2_nand2_1
X_3224_ _2648_ net1044 net842 VPWR VGND sg13g2_nand2_2
X_6012_ net42 VGND VPWR net901 mydesign.accum\[50\] clknet_leaf_23_clk sg13g2_dfrbpq_2
.ends

