module heichips25_systolicArrayTop (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire \mydesign.accum[0] ;
 wire \mydesign.accum[100] ;
 wire \mydesign.accum[101] ;
 wire \mydesign.accum[102] ;
 wire \mydesign.accum[103] ;
 wire \mydesign.accum[104] ;
 wire \mydesign.accum[105] ;
 wire \mydesign.accum[106] ;
 wire \mydesign.accum[107] ;
 wire \mydesign.accum[108] ;
 wire \mydesign.accum[109] ;
 wire \mydesign.accum[10] ;
 wire \mydesign.accum[110] ;
 wire \mydesign.accum[111] ;
 wire \mydesign.accum[112] ;
 wire \mydesign.accum[113] ;
 wire \mydesign.accum[114] ;
 wire \mydesign.accum[115] ;
 wire \mydesign.accum[116] ;
 wire \mydesign.accum[117] ;
 wire \mydesign.accum[118] ;
 wire \mydesign.accum[119] ;
 wire \mydesign.accum[11] ;
 wire \mydesign.accum[120] ;
 wire \mydesign.accum[121] ;
 wire \mydesign.accum[122] ;
 wire \mydesign.accum[123] ;
 wire \mydesign.accum[124] ;
 wire \mydesign.accum[125] ;
 wire \mydesign.accum[126] ;
 wire \mydesign.accum[127] ;
 wire \mydesign.accum[12] ;
 wire \mydesign.accum[13] ;
 wire \mydesign.accum[14] ;
 wire \mydesign.accum[15] ;
 wire \mydesign.accum[16] ;
 wire \mydesign.accum[17] ;
 wire \mydesign.accum[18] ;
 wire \mydesign.accum[19] ;
 wire \mydesign.accum[1] ;
 wire \mydesign.accum[20] ;
 wire \mydesign.accum[21] ;
 wire \mydesign.accum[22] ;
 wire \mydesign.accum[23] ;
 wire \mydesign.accum[24] ;
 wire \mydesign.accum[25] ;
 wire \mydesign.accum[26] ;
 wire \mydesign.accum[27] ;
 wire \mydesign.accum[28] ;
 wire \mydesign.accum[29] ;
 wire \mydesign.accum[2] ;
 wire \mydesign.accum[30] ;
 wire \mydesign.accum[31] ;
 wire \mydesign.accum[32] ;
 wire \mydesign.accum[33] ;
 wire \mydesign.accum[34] ;
 wire \mydesign.accum[35] ;
 wire \mydesign.accum[36] ;
 wire \mydesign.accum[37] ;
 wire \mydesign.accum[38] ;
 wire \mydesign.accum[39] ;
 wire \mydesign.accum[3] ;
 wire \mydesign.accum[40] ;
 wire \mydesign.accum[41] ;
 wire \mydesign.accum[42] ;
 wire \mydesign.accum[43] ;
 wire \mydesign.accum[44] ;
 wire \mydesign.accum[45] ;
 wire \mydesign.accum[46] ;
 wire \mydesign.accum[47] ;
 wire \mydesign.accum[48] ;
 wire \mydesign.accum[49] ;
 wire \mydesign.accum[4] ;
 wire \mydesign.accum[50] ;
 wire \mydesign.accum[51] ;
 wire \mydesign.accum[52] ;
 wire \mydesign.accum[53] ;
 wire \mydesign.accum[54] ;
 wire \mydesign.accum[55] ;
 wire \mydesign.accum[56] ;
 wire \mydesign.accum[57] ;
 wire \mydesign.accum[58] ;
 wire \mydesign.accum[59] ;
 wire \mydesign.accum[5] ;
 wire \mydesign.accum[60] ;
 wire \mydesign.accum[61] ;
 wire \mydesign.accum[62] ;
 wire \mydesign.accum[63] ;
 wire \mydesign.accum[64] ;
 wire \mydesign.accum[65] ;
 wire \mydesign.accum[66] ;
 wire \mydesign.accum[67] ;
 wire \mydesign.accum[68] ;
 wire \mydesign.accum[69] ;
 wire \mydesign.accum[6] ;
 wire \mydesign.accum[70] ;
 wire \mydesign.accum[71] ;
 wire \mydesign.accum[72] ;
 wire \mydesign.accum[73] ;
 wire \mydesign.accum[74] ;
 wire \mydesign.accum[75] ;
 wire \mydesign.accum[76] ;
 wire \mydesign.accum[77] ;
 wire \mydesign.accum[78] ;
 wire \mydesign.accum[79] ;
 wire \mydesign.accum[7] ;
 wire \mydesign.accum[80] ;
 wire \mydesign.accum[81] ;
 wire \mydesign.accum[82] ;
 wire \mydesign.accum[83] ;
 wire \mydesign.accum[84] ;
 wire \mydesign.accum[85] ;
 wire \mydesign.accum[86] ;
 wire \mydesign.accum[87] ;
 wire \mydesign.accum[88] ;
 wire \mydesign.accum[89] ;
 wire \mydesign.accum[8] ;
 wire \mydesign.accum[90] ;
 wire \mydesign.accum[91] ;
 wire \mydesign.accum[92] ;
 wire \mydesign.accum[93] ;
 wire \mydesign.accum[94] ;
 wire \mydesign.accum[95] ;
 wire \mydesign.accum[96] ;
 wire \mydesign.accum[97] ;
 wire \mydesign.accum[98] ;
 wire \mydesign.accum[99] ;
 wire \mydesign.accum[9] ;
 wire \mydesign.compute_en ;
 wire \mydesign.cp2[0] ;
 wire \mydesign.cp2[1] ;
 wire \mydesign.cp2[2] ;
 wire \mydesign.cp[0] ;
 wire \mydesign.cp[1] ;
 wire \mydesign.cp[2] ;
 wire \mydesign.inputs[0][12] ;
 wire \mydesign.inputs[0][13] ;
 wire \mydesign.inputs[0][14] ;
 wire \mydesign.inputs[0][15] ;
 wire \mydesign.inputs[0][16] ;
 wire \mydesign.inputs[0][17] ;
 wire \mydesign.inputs[0][18] ;
 wire \mydesign.inputs[0][19] ;
 wire \mydesign.inputs[0][20] ;
 wire \mydesign.inputs[0][21] ;
 wire \mydesign.inputs[0][22] ;
 wire \mydesign.inputs[0][23] ;
 wire \mydesign.inputs[0][24] ;
 wire \mydesign.inputs[0][25] ;
 wire \mydesign.inputs[0][26] ;
 wire \mydesign.inputs[0][27] ;
 wire \mydesign.inputs[1][10] ;
 wire \mydesign.inputs[1][11] ;
 wire \mydesign.inputs[1][12] ;
 wire \mydesign.inputs[1][13] ;
 wire \mydesign.inputs[1][14] ;
 wire \mydesign.inputs[1][15] ;
 wire \mydesign.inputs[1][16] ;
 wire \mydesign.inputs[1][17] ;
 wire \mydesign.inputs[1][18] ;
 wire \mydesign.inputs[1][19] ;
 wire \mydesign.inputs[1][20] ;
 wire \mydesign.inputs[1][21] ;
 wire \mydesign.inputs[1][22] ;
 wire \mydesign.inputs[1][23] ;
 wire \mydesign.inputs[1][8] ;
 wire \mydesign.inputs[1][9] ;
 wire \mydesign.inputs[2][10] ;
 wire \mydesign.inputs[2][11] ;
 wire \mydesign.inputs[2][12] ;
 wire \mydesign.inputs[2][13] ;
 wire \mydesign.inputs[2][14] ;
 wire \mydesign.inputs[2][15] ;
 wire \mydesign.inputs[2][16] ;
 wire \mydesign.inputs[2][17] ;
 wire \mydesign.inputs[2][18] ;
 wire \mydesign.inputs[2][19] ;
 wire \mydesign.inputs[2][4] ;
 wire \mydesign.inputs[2][5] ;
 wire \mydesign.inputs[2][6] ;
 wire \mydesign.inputs[2][7] ;
 wire \mydesign.inputs[2][8] ;
 wire \mydesign.inputs[2][9] ;
 wire \mydesign.inputs[3][0] ;
 wire \mydesign.inputs[3][10] ;
 wire \mydesign.inputs[3][11] ;
 wire \mydesign.inputs[3][12] ;
 wire \mydesign.inputs[3][13] ;
 wire \mydesign.inputs[3][14] ;
 wire \mydesign.inputs[3][15] ;
 wire \mydesign.inputs[3][1] ;
 wire \mydesign.inputs[3][2] ;
 wire \mydesign.inputs[3][3] ;
 wire \mydesign.inputs[3][4] ;
 wire \mydesign.inputs[3][5] ;
 wire \mydesign.inputs[3][6] ;
 wire \mydesign.inputs[3][7] ;
 wire \mydesign.inputs[3][8] ;
 wire \mydesign.inputs[3][9] ;
 wire \mydesign.load_counter[0] ;
 wire \mydesign.load_counter[1] ;
 wire \mydesign.load_counter[2] ;
 wire \mydesign.load_counter[3] ;
 wire \mydesign.out[0] ;
 wire \mydesign.out[1] ;
 wire \mydesign.out[2] ;
 wire \mydesign.out[3] ;
 wire \mydesign.pe_inputs[10] ;
 wire \mydesign.pe_inputs[11] ;
 wire \mydesign.pe_inputs[12] ;
 wire \mydesign.pe_inputs[13] ;
 wire \mydesign.pe_inputs[14] ;
 wire \mydesign.pe_inputs[15] ;
 wire \mydesign.pe_inputs[20] ;
 wire \mydesign.pe_inputs[21] ;
 wire \mydesign.pe_inputs[22] ;
 wire \mydesign.pe_inputs[23] ;
 wire \mydesign.pe_inputs[24] ;
 wire \mydesign.pe_inputs[25] ;
 wire \mydesign.pe_inputs[26] ;
 wire \mydesign.pe_inputs[27] ;
 wire \mydesign.pe_inputs[28] ;
 wire \mydesign.pe_inputs[29] ;
 wire \mydesign.pe_inputs[30] ;
 wire \mydesign.pe_inputs[31] ;
 wire \mydesign.pe_inputs[36] ;
 wire \mydesign.pe_inputs[37] ;
 wire \mydesign.pe_inputs[38] ;
 wire \mydesign.pe_inputs[39] ;
 wire \mydesign.pe_inputs[40] ;
 wire \mydesign.pe_inputs[41] ;
 wire \mydesign.pe_inputs[42] ;
 wire \mydesign.pe_inputs[43] ;
 wire \mydesign.pe_inputs[44] ;
 wire \mydesign.pe_inputs[45] ;
 wire \mydesign.pe_inputs[46] ;
 wire \mydesign.pe_inputs[47] ;
 wire \mydesign.pe_inputs[4] ;
 wire \mydesign.pe_inputs[52] ;
 wire \mydesign.pe_inputs[53] ;
 wire \mydesign.pe_inputs[54] ;
 wire \mydesign.pe_inputs[55] ;
 wire \mydesign.pe_inputs[56] ;
 wire \mydesign.pe_inputs[57] ;
 wire \mydesign.pe_inputs[58] ;
 wire \mydesign.pe_inputs[59] ;
 wire \mydesign.pe_inputs[5] ;
 wire \mydesign.pe_inputs[60] ;
 wire \mydesign.pe_inputs[61] ;
 wire \mydesign.pe_inputs[62] ;
 wire \mydesign.pe_inputs[63] ;
 wire \mydesign.pe_inputs[6] ;
 wire \mydesign.pe_inputs[7] ;
 wire \mydesign.pe_inputs[8] ;
 wire \mydesign.pe_inputs[9] ;
 wire \mydesign.pe_weights[16] ;
 wire \mydesign.pe_weights[17] ;
 wire \mydesign.pe_weights[18] ;
 wire \mydesign.pe_weights[19] ;
 wire \mydesign.pe_weights[20] ;
 wire \mydesign.pe_weights[21] ;
 wire \mydesign.pe_weights[22] ;
 wire \mydesign.pe_weights[23] ;
 wire \mydesign.pe_weights[24] ;
 wire \mydesign.pe_weights[25] ;
 wire \mydesign.pe_weights[26] ;
 wire \mydesign.pe_weights[27] ;
 wire \mydesign.pe_weights[28] ;
 wire \mydesign.pe_weights[29] ;
 wire \mydesign.pe_weights[30] ;
 wire \mydesign.pe_weights[31] ;
 wire \mydesign.pe_weights[32] ;
 wire \mydesign.pe_weights[33] ;
 wire \mydesign.pe_weights[34] ;
 wire \mydesign.pe_weights[35] ;
 wire \mydesign.pe_weights[36] ;
 wire \mydesign.pe_weights[37] ;
 wire \mydesign.pe_weights[38] ;
 wire \mydesign.pe_weights[39] ;
 wire \mydesign.pe_weights[40] ;
 wire \mydesign.pe_weights[41] ;
 wire \mydesign.pe_weights[42] ;
 wire \mydesign.pe_weights[43] ;
 wire \mydesign.pe_weights[44] ;
 wire \mydesign.pe_weights[45] ;
 wire \mydesign.pe_weights[46] ;
 wire \mydesign.pe_weights[47] ;
 wire \mydesign.pe_weights[48] ;
 wire \mydesign.pe_weights[49] ;
 wire \mydesign.pe_weights[50] ;
 wire \mydesign.pe_weights[51] ;
 wire \mydesign.pe_weights[52] ;
 wire \mydesign.pe_weights[53] ;
 wire \mydesign.pe_weights[54] ;
 wire \mydesign.pe_weights[55] ;
 wire \mydesign.pe_weights[56] ;
 wire \mydesign.pe_weights[57] ;
 wire \mydesign.pe_weights[58] ;
 wire \mydesign.pe_weights[59] ;
 wire \mydesign.pe_weights[60] ;
 wire \mydesign.pe_weights[61] ;
 wire \mydesign.pe_weights[62] ;
 wire \mydesign.pe_weights[63] ;
 wire \mydesign.valid_out ;
 wire \mydesign.weights[0][12] ;
 wire \mydesign.weights[0][13] ;
 wire \mydesign.weights[0][14] ;
 wire \mydesign.weights[0][15] ;
 wire \mydesign.weights[0][16] ;
 wire \mydesign.weights[0][17] ;
 wire \mydesign.weights[0][18] ;
 wire \mydesign.weights[0][19] ;
 wire \mydesign.weights[0][20] ;
 wire \mydesign.weights[0][21] ;
 wire \mydesign.weights[0][22] ;
 wire \mydesign.weights[0][23] ;
 wire \mydesign.weights[0][24] ;
 wire \mydesign.weights[0][25] ;
 wire \mydesign.weights[0][26] ;
 wire \mydesign.weights[0][27] ;
 wire \mydesign.weights[1][10] ;
 wire \mydesign.weights[1][11] ;
 wire \mydesign.weights[1][12] ;
 wire \mydesign.weights[1][13] ;
 wire \mydesign.weights[1][14] ;
 wire \mydesign.weights[1][15] ;
 wire \mydesign.weights[1][16] ;
 wire \mydesign.weights[1][17] ;
 wire \mydesign.weights[1][18] ;
 wire \mydesign.weights[1][19] ;
 wire \mydesign.weights[1][20] ;
 wire \mydesign.weights[1][21] ;
 wire \mydesign.weights[1][22] ;
 wire \mydesign.weights[1][23] ;
 wire \mydesign.weights[1][8] ;
 wire \mydesign.weights[1][9] ;
 wire \mydesign.weights[2][10] ;
 wire \mydesign.weights[2][11] ;
 wire \mydesign.weights[2][12] ;
 wire \mydesign.weights[2][13] ;
 wire \mydesign.weights[2][14] ;
 wire \mydesign.weights[2][15] ;
 wire \mydesign.weights[2][16] ;
 wire \mydesign.weights[2][17] ;
 wire \mydesign.weights[2][18] ;
 wire \mydesign.weights[2][19] ;
 wire \mydesign.weights[2][4] ;
 wire \mydesign.weights[2][5] ;
 wire \mydesign.weights[2][6] ;
 wire \mydesign.weights[2][7] ;
 wire \mydesign.weights[2][8] ;
 wire \mydesign.weights[2][9] ;
 wire \mydesign.weights[3][0] ;
 wire \mydesign.weights[3][10] ;
 wire \mydesign.weights[3][11] ;
 wire \mydesign.weights[3][12] ;
 wire \mydesign.weights[3][13] ;
 wire \mydesign.weights[3][14] ;
 wire \mydesign.weights[3][15] ;
 wire \mydesign.weights[3][1] ;
 wire \mydesign.weights[3][2] ;
 wire \mydesign.weights[3][3] ;
 wire \mydesign.weights[3][4] ;
 wire \mydesign.weights[3][5] ;
 wire \mydesign.weights[3][6] ;
 wire \mydesign.weights[3][7] ;
 wire \mydesign.weights[3][8] ;
 wire \mydesign.weights[3][9] ;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire clknet_leaf_0_clk;
 wire net7;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net16;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;

 sg13g2_inv_4 _3075_ (.A(net590),
    .Y(_2516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3076_ (.Y(_2517_),
    .A(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3077_ (.Y(_2518_),
    .A(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3078_ (.Y(_2519_),
    .A(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3079_ (.Y(_2520_),
    .A(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3080_ (.VDD(VPWR),
    .Y(_2521_),
    .A(net520),
    .VSS(VGND));
 sg13g2_inv_1 _3081_ (.VDD(VPWR),
    .Y(_2522_),
    .A(net832),
    .VSS(VGND));
 sg13g2_inv_1 _3082_ (.VDD(VPWR),
    .Y(_2523_),
    .A(net934),
    .VSS(VGND));
 sg13g2_inv_1 _3083_ (.VDD(VPWR),
    .Y(_2524_),
    .A(net521),
    .VSS(VGND));
 sg13g2_inv_1 _3084_ (.VDD(VPWR),
    .Y(_2525_),
    .A(net1000),
    .VSS(VGND));
 sg13g2_inv_1 _3085_ (.VDD(VPWR),
    .Y(_2526_),
    .A(net939),
    .VSS(VGND));
 sg13g2_inv_1 _3086_ (.VDD(VPWR),
    .Y(_2527_),
    .A(net522),
    .VSS(VGND));
 sg13g2_inv_1 _3087_ (.VDD(VPWR),
    .Y(_2528_),
    .A(net773),
    .VSS(VGND));
 sg13g2_inv_1 _3088_ (.VDD(VPWR),
    .Y(_2529_),
    .A(net816),
    .VSS(VGND));
 sg13g2_inv_1 _3089_ (.VDD(VPWR),
    .Y(_2530_),
    .A(net530),
    .VSS(VGND));
 sg13g2_inv_1 _3090_ (.VDD(VPWR),
    .Y(_2531_),
    .A(net828),
    .VSS(VGND));
 sg13g2_inv_1 _3091_ (.VDD(VPWR),
    .Y(_2532_),
    .A(net1033),
    .VSS(VGND));
 sg13g2_inv_1 _3092_ (.VDD(VPWR),
    .Y(_2533_),
    .A(net531),
    .VSS(VGND));
 sg13g2_inv_1 _3093_ (.VDD(VPWR),
    .Y(_2534_),
    .A(net830),
    .VSS(VGND));
 sg13g2_inv_1 _3094_ (.VDD(VPWR),
    .Y(_2535_),
    .A(net862),
    .VSS(VGND));
 sg13g2_inv_1 _3095_ (.VDD(VPWR),
    .Y(_2536_),
    .A(net943),
    .VSS(VGND));
 sg13g2_inv_1 _3096_ (.VDD(VPWR),
    .Y(_2537_),
    .A(net974),
    .VSS(VGND));
 sg13g2_inv_1 _3097_ (.VDD(VPWR),
    .Y(_2538_),
    .A(net1031),
    .VSS(VGND));
 sg13g2_inv_1 _3098_ (.VDD(VPWR),
    .Y(_2539_),
    .A(net849),
    .VSS(VGND));
 sg13g2_inv_1 _3099_ (.VDD(VPWR),
    .Y(_2540_),
    .A(net528),
    .VSS(VGND));
 sg13g2_inv_1 _3100_ (.VDD(VPWR),
    .Y(_2541_),
    .A(net789),
    .VSS(VGND));
 sg13g2_inv_1 _3101_ (.VDD(VPWR),
    .Y(_2542_),
    .A(net813),
    .VSS(VGND));
 sg13g2_inv_1 _3102_ (.VDD(VPWR),
    .Y(_2543_),
    .A(net856),
    .VSS(VGND));
 sg13g2_inv_1 _3103_ (.VDD(VPWR),
    .Y(_2544_),
    .A(net1013),
    .VSS(VGND));
 sg13g2_inv_1 _3104_ (.VDD(VPWR),
    .Y(_2545_),
    .A(net887),
    .VSS(VGND));
 sg13g2_inv_1 _3105_ (.VDD(VPWR),
    .Y(_2546_),
    .A(net879),
    .VSS(VGND));
 sg13g2_inv_2 _3106_ (.Y(_2547_),
    .A(net529),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3107_ (.VDD(VPWR),
    .Y(_2548_),
    .A(\mydesign.accum[61] ),
    .VSS(VGND));
 sg13g2_inv_1 _3108_ (.VDD(VPWR),
    .Y(_2549_),
    .A(net535),
    .VSS(VGND));
 sg13g2_inv_1 _3109_ (.VDD(VPWR),
    .Y(_2550_),
    .A(net952),
    .VSS(VGND));
 sg13g2_inv_1 _3110_ (.VDD(VPWR),
    .Y(_2551_),
    .A(net811),
    .VSS(VGND));
 sg13g2_inv_1 _3111_ (.VDD(VPWR),
    .Y(_2552_),
    .A(net815),
    .VSS(VGND));
 sg13g2_inv_2 _3112_ (.Y(_2553_),
    .A(net537),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3113_ (.Y(_2554_),
    .A(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3114_ (.Y(_2555_),
    .A(net872),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3115_ (.VDD(VPWR),
    .Y(_2556_),
    .A(net538),
    .VSS(VGND));
 sg13g2_inv_1 _3116_ (.VDD(VPWR),
    .Y(_2557_),
    .A(net996),
    .VSS(VGND));
 sg13g2_inv_1 _3117_ (.VDD(VPWR),
    .Y(_2558_),
    .A(net971),
    .VSS(VGND));
 sg13g2_inv_2 _3118_ (.Y(_2559_),
    .A(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3119_ (.VDD(VPWR),
    .Y(_2560_),
    .A(net993),
    .VSS(VGND));
 sg13g2_inv_1 _3120_ (.VDD(VPWR),
    .Y(_2561_),
    .A(net981),
    .VSS(VGND));
 sg13g2_inv_1 _3121_ (.VDD(VPWR),
    .Y(_2562_),
    .A(net899),
    .VSS(VGND));
 sg13g2_inv_1 _3122_ (.VDD(VPWR),
    .Y(_2563_),
    .A(net534),
    .VSS(VGND));
 sg13g2_inv_1 _3123_ (.VDD(VPWR),
    .Y(_2564_),
    .A(net539),
    .VSS(VGND));
 sg13g2_inv_1 _3124_ (.VDD(VPWR),
    .Y(_2565_),
    .A(net988),
    .VSS(VGND));
 sg13g2_inv_1 _3125_ (.VDD(VPWR),
    .Y(_2566_),
    .A(net989),
    .VSS(VGND));
 sg13g2_inv_2 _3126_ (.Y(_2567_),
    .A(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3127_ (.Y(_2568_),
    .A(net956),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3128_ (.VDD(VPWR),
    .Y(_2569_),
    .A(net1082),
    .VSS(VGND));
 sg13g2_inv_2 _3129_ (.Y(_2570_),
    .A(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3130_ (.Y(_2571_),
    .A(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3131_ (.VDD(VPWR),
    .Y(_2572_),
    .A(\mydesign.accum[94] ),
    .VSS(VGND));
 sg13g2_inv_1 _3132_ (.VDD(VPWR),
    .Y(_2573_),
    .A(net999),
    .VSS(VGND));
 sg13g2_inv_1 _3133_ (.VDD(VPWR),
    .Y(_2574_),
    .A(net804),
    .VSS(VGND));
 sg13g2_inv_1 _3134_ (.VDD(VPWR),
    .Y(_2575_),
    .A(net881),
    .VSS(VGND));
 sg13g2_inv_1 _3135_ (.VDD(VPWR),
    .Y(_2576_),
    .A(net838),
    .VSS(VGND));
 sg13g2_inv_1 _3136_ (.VDD(VPWR),
    .Y(_2577_),
    .A(net880),
    .VSS(VGND));
 sg13g2_inv_1 _3137_ (.VDD(VPWR),
    .Y(_2578_),
    .A(net808),
    .VSS(VGND));
 sg13g2_inv_1 _3138_ (.VDD(VPWR),
    .Y(_2579_),
    .A(net757),
    .VSS(VGND));
 sg13g2_inv_1 _3139_ (.VDD(VPWR),
    .Y(_2580_),
    .A(net1046),
    .VSS(VGND));
 sg13g2_inv_1 _3140_ (.VDD(VPWR),
    .Y(_2581_),
    .A(net1027),
    .VSS(VGND));
 sg13g2_inv_1 _3141_ (.VDD(VPWR),
    .Y(_2582_),
    .A(net1015),
    .VSS(VGND));
 sg13g2_inv_1 _3142_ (.VDD(VPWR),
    .Y(_2583_),
    .A(net1073),
    .VSS(VGND));
 sg13g2_inv_1 _3143_ (.VDD(VPWR),
    .Y(_2584_),
    .A(net407),
    .VSS(VGND));
 sg13g2_inv_1 _3144_ (.VDD(VPWR),
    .Y(_2585_),
    .A(net756),
    .VSS(VGND));
 sg13g2_inv_4 _3145_ (.A(net541),
    .Y(_2586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3146_ (.Y(_2587_),
    .A(net547),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3147_ (.Y(_2588_),
    .A(net1110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3148_ (.VDD(VPWR),
    .Y(_2589_),
    .A(\mydesign.weights[2][16] ),
    .VSS(VGND));
 sg13g2_inv_1 _3149_ (.VDD(VPWR),
    .Y(_2590_),
    .A(net623),
    .VSS(VGND));
 sg13g2_inv_8 _3150_ (.Y(_2591_),
    .A(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3151_ (.VDD(VPWR),
    .Y(_2592_),
    .A(\mydesign.weights[0][24] ),
    .VSS(VGND));
 sg13g2_inv_1 _3152_ (.VDD(VPWR),
    .Y(_2593_),
    .A(net411),
    .VSS(VGND));
 sg13g2_inv_1 _3153_ (.VDD(VPWR),
    .Y(_2594_),
    .A(\mydesign.inputs[2][7] ),
    .VSS(VGND));
 sg13g2_nor2b_2 _3154_ (.A(net555),
    .B_N(net545),
    .Y(_2595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3155_ (.A(net541),
    .B(net496),
    .X(_2596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3156_ (.Y(_2597_),
    .A(net541),
    .B(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3157_ (.B(net756),
    .C(net744),
    .A(_2584_),
    .Y(_2598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3158_ (.A(net610),
    .B(net5),
    .Y(_2599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3159_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2600_),
    .B(net5),
    .A(net610));
 sg13g2_nor2_1 _3160_ (.A(net499),
    .B(net611),
    .Y(_2601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3161_ (.Y(_2602_),
    .A(net563),
    .B(_2591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3162_ (.A(net499),
    .B(_2600_),
    .Y(_2603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3163_ (.VDD(VPWR),
    .Y(_2604_),
    .A(_2603_),
    .VSS(VGND));
 sg13g2_nor4_1 _3164_ (.A(net607),
    .B(_2597_),
    .C(_2598_),
    .D(_2604_),
    .Y(_0000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3165_ (.Y(_2605_),
    .A(net614),
    .B(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3166_ (.Y(_2606_),
    .B(net1106),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\mydesign.load_counter[0] ));
 sg13g2_nand2_2 _3167_ (.Y(_2607_),
    .A(\mydesign.load_counter[3] ),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3168_ (.A(_2605_),
    .B(_2606_),
    .C(_2607_),
    .Y(_2608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3169_ (.Y(_2609_),
    .A(net1),
    .B(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3170_ (.Y(_2610_),
    .A(net747),
    .B(net618),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3171_ (.B1(_2609_),
    .VDD(VPWR),
    .Y(_0001_),
    .VSS(VGND),
    .A1(net432),
    .A2(_2610_));
 sg13g2_nand2_1 _3172_ (.Y(_2611_),
    .A(net2),
    .B(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3173_ (.Y(_2612_),
    .A(net733),
    .B(net616),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3174_ (.B1(_2611_),
    .VDD(VPWR),
    .Y(_0002_),
    .VSS(VGND),
    .A1(net432),
    .A2(_2612_));
 sg13g2_nand2_1 _3175_ (.Y(_2613_),
    .A(net3),
    .B(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3176_ (.Y(_2614_),
    .A(net741),
    .B(net616),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3177_ (.B1(_2613_),
    .VDD(VPWR),
    .Y(_0003_),
    .VSS(VGND),
    .A1(net432),
    .A2(_2614_));
 sg13g2_nand2_1 _3178_ (.Y(_2615_),
    .A(net4),
    .B(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3179_ (.Y(_2616_),
    .A(net752),
    .B(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3180_ (.B1(_2615_),
    .VDD(VPWR),
    .Y(_0004_),
    .VSS(VGND),
    .A1(_2608_),
    .A2(_2616_));
 sg13g2_nor2b_2 _3181_ (.A(net610),
    .B_N(net5),
    .Y(_2617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3182_ (.Y(_2618_),
    .A(_2591_),
    .B(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3183_ (.A(net1044),
    .B(net842),
    .Y(_2619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3184_ (.VDD(VPWR),
    .Y(_2620_),
    .A(_2619_),
    .VSS(VGND));
 sg13g2_nor2_1 _3185_ (.A(\mydesign.load_counter[3] ),
    .B(net596),
    .Y(_2621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3186_ (.Y(_2622_),
    .A(_2621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3187_ (.B(_2619_),
    .C(_2621_),
    .A(net605),
    .Y(_2623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3188_ (.B(net754),
    .C(_2623_),
    .A(net620),
    .Y(_2624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3189_ (.Y(_2625_),
    .A(net1),
    .B(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3190_ (.B1(_2624_),
    .VDD(VPWR),
    .Y(_0005_),
    .VSS(VGND),
    .A1(_2623_),
    .A2(net603));
 sg13g2_nand3_1 _3191_ (.B(net760),
    .C(_2623_),
    .A(net621),
    .Y(_2626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3192_ (.Y(_2627_),
    .A(net2),
    .B(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3193_ (.B1(_2626_),
    .VDD(VPWR),
    .Y(_0006_),
    .VSS(VGND),
    .A1(_2623_),
    .A2(net601));
 sg13g2_nand3_1 _3194_ (.B(net728),
    .C(_2623_),
    .A(net620),
    .Y(_2628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3195_ (.Y(_2629_),
    .A(net3),
    .B(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3196_ (.B1(_2628_),
    .VDD(VPWR),
    .Y(_0007_),
    .VSS(VGND),
    .A1(_2623_),
    .A2(net600));
 sg13g2_nand3_1 _3197_ (.B(net738),
    .C(_2623_),
    .A(net620),
    .Y(_2630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3198_ (.Y(_2631_),
    .A(net4),
    .B(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3199_ (.B1(_2630_),
    .VDD(VPWR),
    .Y(_0008_),
    .VSS(VGND),
    .A1(_2623_),
    .A2(net598));
 sg13g2_nor2_2 _3200_ (.A(_2606_),
    .B(_2622_),
    .Y(_2632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3201_ (.Y(_2633_),
    .B(_2632_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2605_));
 sg13g2_nand3_1 _3202_ (.B(net617),
    .C(_2633_),
    .A(net677),
    .Y(_2634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3203_ (.B1(_2634_),
    .VDD(VPWR),
    .Y(_0009_),
    .VSS(VGND),
    .A1(_2520_),
    .A2(_2633_));
 sg13g2_nand3_1 _3204_ (.B(net616),
    .C(_2633_),
    .A(net675),
    .Y(_2635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3205_ (.B1(_2635_),
    .VDD(VPWR),
    .Y(_0010_),
    .VSS(VGND),
    .A1(_2519_),
    .A2(_2633_));
 sg13g2_nand3_1 _3206_ (.B(net616),
    .C(_2633_),
    .A(net692),
    .Y(_2636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3207_ (.B1(_2636_),
    .VDD(VPWR),
    .Y(_0011_),
    .VSS(VGND),
    .A1(_2518_),
    .A2(_2633_));
 sg13g2_nand3_1 _3208_ (.B(net617),
    .C(_2633_),
    .A(net662),
    .Y(_2637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3209_ (.B1(_2637_),
    .VDD(VPWR),
    .Y(_0012_),
    .VSS(VGND),
    .A1(_2517_),
    .A2(_2633_));
 sg13g2_nor2_1 _3210_ (.A(_2588_),
    .B(net596),
    .Y(_2638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3211_ (.Y(_2639_),
    .B(\mydesign.load_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1108));
 sg13g2_nor2_2 _3212_ (.A(_2606_),
    .B(_2639_),
    .Y(_2640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3213_ (.Y(_2641_),
    .A(net606),
    .B(_2640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3214_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net609),
    .Y(_2642_),
    .A2(_2640_),
    .A1(net605));
 sg13g2_nand2_1 _3215_ (.Y(_2643_),
    .A(net423),
    .B(_2642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3216_ (.B1(_2643_),
    .VDD(VPWR),
    .Y(_0013_),
    .VSS(VGND),
    .A1(net604),
    .A2(_2641_));
 sg13g2_nand2_1 _3217_ (.Y(_2644_),
    .A(net420),
    .B(_2642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3218_ (.B1(_2644_),
    .VDD(VPWR),
    .Y(_0014_),
    .VSS(VGND),
    .A1(net602),
    .A2(_2641_));
 sg13g2_nand2_1 _3219_ (.Y(_2645_),
    .A(net667),
    .B(_2642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3220_ (.B1(_2645_),
    .VDD(VPWR),
    .Y(_0015_),
    .VSS(VGND),
    .A1(net600),
    .A2(_2641_));
 sg13g2_nand2_1 _3221_ (.Y(_2646_),
    .A(net642),
    .B(_2642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3222_ (.B1(_2646_),
    .VDD(VPWR),
    .Y(_0016_),
    .VSS(VGND),
    .A1(net598),
    .A2(_2641_));
 sg13g2_and2_1 _3223_ (.A(net1044),
    .B(net842),
    .X(_2647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3224_ (.Y(_2648_),
    .A(net1044),
    .B(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3225_ (.B(_2638_),
    .C(_2647_),
    .A(net605),
    .Y(_2649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3226_ (.A(net623),
    .B(_2649_),
    .X(_2650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3227_ (.Y(_2651_),
    .A(net655),
    .B(_2650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3228_ (.B1(_2651_),
    .VDD(VPWR),
    .Y(_0017_),
    .VSS(VGND),
    .A1(net604),
    .A2(_2649_));
 sg13g2_nand2_1 _3229_ (.Y(_2652_),
    .A(net413),
    .B(_2650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3230_ (.B1(_2652_),
    .VDD(VPWR),
    .Y(_0018_),
    .VSS(VGND),
    .A1(net602),
    .A2(_2649_));
 sg13g2_nand2_1 _3231_ (.Y(_2653_),
    .A(net704),
    .B(_2650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3232_ (.B1(_2653_),
    .VDD(VPWR),
    .Y(_0019_),
    .VSS(VGND),
    .A1(net600),
    .A2(_2649_));
 sg13g2_nand2_1 _3233_ (.Y(_2654_),
    .A(net669),
    .B(_2650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3234_ (.B1(_2654_),
    .VDD(VPWR),
    .Y(_0020_),
    .VSS(VGND),
    .A1(net598),
    .A2(_2649_));
 sg13g2_nand2_2 _3235_ (.Y(_2655_),
    .A(net614),
    .B(_2618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3236_ (.A(net596),
    .B(_2647_),
    .X(_2656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3237_ (.Y(_2657_),
    .A(_2588_),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3238_ (.A(_2648_),
    .B(_2657_),
    .Y(_2658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _3239_ (.A2(_2658_),
    .A1(net605),
    .B1(net607),
    .X(_2659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3240_ (.A(net608),
    .B(net611),
    .Y(_2660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3241_ (.Y(_2661_),
    .A(net617),
    .B(_2591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3242_ (.Y(_2662_),
    .A(net614),
    .B(net605),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3243_ (.A(_2620_),
    .B(net1109),
    .Y(_2663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3244_ (.A(_2632_),
    .B(_2663_),
    .Y(_2664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3245_ (.B1(_2588_),
    .VDD(VPWR),
    .Y(_2665_),
    .VSS(VGND),
    .A1(net596),
    .A2(\mydesign.load_counter[0] ));
 sg13g2_a21oi_2 _3246_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2662_),
    .Y(_2666_),
    .A2(_2665_),
    .A1(_2664_));
 sg13g2_and2_1 _3247_ (.A(net1),
    .B(_2666_),
    .X(_2667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3248_ (.A0(net794),
    .A1(_2667_),
    .S(_2659_),
    .X(_0021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3249_ (.A(net2),
    .B(_2666_),
    .X(_2668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3250_ (.A0(net799),
    .A1(_2668_),
    .S(_2659_),
    .X(_0022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3251_ (.A(net3),
    .B(_2666_),
    .X(_2669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3252_ (.A0(net791),
    .A1(_2669_),
    .S(_2659_),
    .X(_0023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3253_ (.A(net4),
    .B(_2666_),
    .X(_2670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3254_ (.A0(net800),
    .A1(_2670_),
    .S(_2659_),
    .X(_0024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3255_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2671_),
    .B(_2657_),
    .A(_2606_));
 sg13g2_o21ai_1 _3256_ (.B1(net614),
    .VDD(VPWR),
    .Y(_2672_),
    .VSS(VGND),
    .A1(_2618_),
    .A2(_2671_));
 sg13g2_mux2_1 _3257_ (.A0(net762),
    .A1(_2667_),
    .S(_2672_),
    .X(_0025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3258_ (.A0(net769),
    .A1(_2668_),
    .S(_2672_),
    .X(_0026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3259_ (.A0(net797),
    .A1(_2669_),
    .S(_2672_),
    .X(_0027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3260_ (.A0(net775),
    .A1(_2670_),
    .S(_2672_),
    .X(_0028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3261_ (.A(_2591_),
    .B(_2671_),
    .Y(_2673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3262_ (.B1(net617),
    .VDD(VPWR),
    .Y(_2674_),
    .VSS(VGND),
    .A1(net805),
    .A2(_2673_));
 sg13g2_a21oi_1 _3263_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2520_),
    .A2(_2673_),
    .Y(_0029_),
    .B1(_2674_));
 sg13g2_o21ai_1 _3264_ (.B1(net616),
    .VDD(VPWR),
    .Y(_2675_),
    .VSS(VGND),
    .A1(net807),
    .A2(_2673_));
 sg13g2_a21oi_1 _3265_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2519_),
    .A2(_2673_),
    .Y(_0030_),
    .B1(_2675_));
 sg13g2_o21ai_1 _3266_ (.B1(net616),
    .VDD(VPWR),
    .Y(_2676_),
    .VSS(VGND),
    .A1(net810),
    .A2(_2673_));
 sg13g2_a21oi_1 _3267_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2518_),
    .A2(_2673_),
    .Y(_0031_),
    .B1(_2676_));
 sg13g2_o21ai_1 _3268_ (.B1(net617),
    .VDD(VPWR),
    .Y(_2677_),
    .VSS(VGND),
    .A1(net885),
    .A2(_2673_));
 sg13g2_a21oi_1 _3269_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2517_),
    .A2(_2673_),
    .Y(_0032_),
    .B1(_2677_));
 sg13g2_nand2b_2 _3270_ (.Y(_2678_),
    .B(_2663_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2662_));
 sg13g2_nand3_1 _3271_ (.B(net617),
    .C(_2678_),
    .A(net670),
    .Y(_2679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3272_ (.B1(_2679_),
    .VDD(VPWR),
    .Y(_0033_),
    .VSS(VGND),
    .A1(_2520_),
    .A2(_2678_));
 sg13g2_nand3_1 _3273_ (.B(net617),
    .C(_2678_),
    .A(net682),
    .Y(_2680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3274_ (.B1(_2680_),
    .VDD(VPWR),
    .Y(_0034_),
    .VSS(VGND),
    .A1(_2519_),
    .A2(_2678_));
 sg13g2_nand3_1 _3275_ (.B(net616),
    .C(_2678_),
    .A(net703),
    .Y(_2681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3276_ (.B1(_2681_),
    .VDD(VPWR),
    .Y(_0035_),
    .VSS(VGND),
    .A1(_2518_),
    .A2(_2678_));
 sg13g2_nand3_1 _3277_ (.B(net616),
    .C(_2678_),
    .A(net736),
    .Y(_2682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3278_ (.B1(_2682_),
    .VDD(VPWR),
    .Y(_0036_),
    .VSS(VGND),
    .A1(_2517_),
    .A2(_2678_));
 sg13g2_nand2b_2 _3279_ (.Y(_2683_),
    .B(\mydesign.load_counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\mydesign.load_counter[1] ));
 sg13g2_o21ai_1 _3280_ (.B1(net614),
    .VDD(VPWR),
    .Y(_2684_),
    .VSS(VGND),
    .A1(_2657_),
    .A2(_2683_));
 sg13g2_nand2_2 _3281_ (.Y(_2685_),
    .A(_2655_),
    .B(_2684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3282_ (.A0(_2667_),
    .A1(net796),
    .S(_2685_),
    .X(_0037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3283_ (.A0(_2668_),
    .A1(net782),
    .S(_2685_),
    .X(_0038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3284_ (.A0(_2669_),
    .A1(net776),
    .S(_2685_),
    .X(_0039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3285_ (.A0(_2670_),
    .A1(net778),
    .S(_2685_),
    .X(_0040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3286_ (.B1(net614),
    .VDD(VPWR),
    .Y(_2686_),
    .VSS(VGND),
    .A1(_2620_),
    .A2(_2657_));
 sg13g2_nand2_2 _3287_ (.Y(_2687_),
    .A(_2655_),
    .B(_2686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3288_ (.A0(_2667_),
    .A1(net795),
    .S(_2687_),
    .X(_0041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3289_ (.A0(_2668_),
    .A1(net779),
    .S(_2687_),
    .X(_0042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3290_ (.A0(_2669_),
    .A1(net793),
    .S(_2687_),
    .X(_0043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3291_ (.A0(_2670_),
    .A1(net798),
    .S(_2687_),
    .X(_0044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3292_ (.Y(_2688_),
    .A(_2588_),
    .B(_2647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3293_ (.A(net596),
    .B(_2688_),
    .Y(_2689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3294_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net608),
    .Y(_2690_),
    .A2(_2689_),
    .A1(net605));
 sg13g2_mux2_1 _3295_ (.A0(_2667_),
    .A1(net765),
    .S(_2690_),
    .X(_0045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3296_ (.A0(_2668_),
    .A1(net786),
    .S(_2690_),
    .X(_0046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3297_ (.A0(_2669_),
    .A1(net772),
    .S(_2690_),
    .X(_0047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3298_ (.A0(_2670_),
    .A1(net787),
    .S(_2690_),
    .X(_0048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _3299_ (.A2(_2632_),
    .A1(net605),
    .B1(net608),
    .X(_2691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3300_ (.A0(net780),
    .A1(_2667_),
    .S(_2691_),
    .X(_0049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3301_ (.A0(net766),
    .A1(_2668_),
    .S(_2691_),
    .X(_0050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3302_ (.A0(net788),
    .A1(_2669_),
    .S(_2691_),
    .X(_0051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3303_ (.A0(net801),
    .A1(_2670_),
    .S(_2691_),
    .X(_0052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3304_ (.B(net605),
    .C(_2656_),
    .A(net1064),
    .Y(_2692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3305_ (.B(net709),
    .C(net429),
    .A(net618),
    .Y(_2693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3306_ (.B1(_2693_),
    .VDD(VPWR),
    .Y(_0053_),
    .VSS(VGND),
    .A1(net603),
    .A2(net429));
 sg13g2_nand3_1 _3307_ (.B(net742),
    .C(net429),
    .A(net618),
    .Y(_2694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3308_ (.B1(_2694_),
    .VDD(VPWR),
    .Y(_0054_),
    .VSS(VGND),
    .A1(net601),
    .A2(net429));
 sg13g2_nand3_1 _3309_ (.B(net712),
    .C(net429),
    .A(net618),
    .Y(_2695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3310_ (.B1(_2695_),
    .VDD(VPWR),
    .Y(_0055_),
    .VSS(VGND),
    .A1(net599),
    .A2(net429));
 sg13g2_nand3_1 _3311_ (.B(net719),
    .C(net429),
    .A(net618),
    .Y(_2696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3312_ (.B1(_2696_),
    .VDD(VPWR),
    .Y(_0056_),
    .VSS(VGND),
    .A1(net597),
    .A2(net429));
 sg13g2_and3_1 _3313_ (.X(_2697_),
    .A(net499),
    .B(net6),
    .C(_2599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3314_ (.B(net6),
    .C(_2599_),
    .A(net499),
    .Y(_2698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3315_ (.A(_2603_),
    .B(net431),
    .Y(_0376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3316_ (.B1(net613),
    .VDD(VPWR),
    .Y(_0377_),
    .VSS(VGND),
    .A1(net842),
    .A2(_2600_));
 sg13g2_a21oi_1 _3317_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net842),
    .A2(_0376_),
    .Y(_0057_),
    .B1(_0377_));
 sg13g2_o21ai_1 _3318_ (.B1(net1044),
    .VDD(VPWR),
    .Y(_0378_),
    .VSS(VGND),
    .A1(_2603_),
    .A2(net431));
 sg13g2_nand3_1 _3319_ (.B(_2620_),
    .C(_2648_),
    .A(_2600_),
    .Y(_0379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3320_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0378_),
    .A2(_0379_),
    .Y(_0058_),
    .B1(net607));
 sg13g2_o21ai_1 _3321_ (.B1(_0376_),
    .VDD(VPWR),
    .Y(_0380_),
    .VSS(VGND),
    .A1(_2599_),
    .A2(_2656_));
 sg13g2_a21oi_1 _3322_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2600_),
    .A2(_2647_),
    .Y(_0381_),
    .B1(net596));
 sg13g2_nand2_1 _3323_ (.Y(_0382_),
    .A(net614),
    .B(_0380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3324_ (.A(_0381_),
    .B(_0382_),
    .Y(_0059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3325_ (.Y(_0383_),
    .B1(_0380_),
    .B2(net1064),
    .A2(_2658_),
    .A1(_2600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3326_ (.A(net607),
    .B(_0383_),
    .Y(_0060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3327_ (.B1(net563),
    .VDD(VPWR),
    .Y(_0384_),
    .VSS(VGND),
    .A1(_2597_),
    .A2(_2598_));
 sg13g2_nand2_1 _3328_ (.Y(_0385_),
    .A(_2692_),
    .B(_0384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3329_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net563),
    .A2(_2600_),
    .Y(_0386_),
    .B1(_0385_));
 sg13g2_nor2_1 _3330_ (.A(net607),
    .B(_0386_),
    .Y(_0061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3331_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2604_),
    .Y(_0387_),
    .A2(_2598_),
    .A1(net454));
 sg13g2_or2_1 _3332_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0388_),
    .B(_0387_),
    .A(net548));
 sg13g2_o21ai_1 _3333_ (.B1(_0387_),
    .VDD(VPWR),
    .Y(_0389_),
    .VSS(VGND),
    .A1(net548),
    .A2(net454));
 sg13g2_and3_1 _3334_ (.X(_0062_),
    .A(net613),
    .B(_0388_),
    .C(_0389_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3335_ (.A(net544),
    .B_N(net555),
    .Y(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3336_ (.Y(_0391_),
    .B1(net461),
    .B2(_0387_),
    .A2(_0389_),
    .A1(net546),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3337_ (.A(net607),
    .B(_0391_),
    .Y(_0063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3338_ (.A(net541),
    .B_N(net546),
    .Y(_0392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3339_ (.Y(_0393_),
    .B(net546),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net543));
 sg13g2_and2_1 _3340_ (.A(net544),
    .B(net554),
    .X(_0394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3341_ (.A(net497),
    .B(_0393_),
    .Y(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3342_ (.A(net545),
    .B_N(net543),
    .Y(_0396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3343_ (.Y(_0397_),
    .B(net541),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net546));
 sg13g2_nor2_1 _3344_ (.A(_0395_),
    .B(net459),
    .Y(_0398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3345_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0398_),
    .C1(net607),
    .B1(_0387_),
    .A1(_2586_),
    .Y(_0064_),
    .A2(_2604_));
 sg13g2_a21oi_1 _3346_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net454),
    .A2(_2603_),
    .Y(_0399_),
    .B1(net744));
 sg13g2_nand4_1 _3347_ (.B(net454),
    .C(_2598_),
    .A(net744),
    .Y(_0400_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2603_));
 sg13g2_nand2_1 _3348_ (.Y(_0401_),
    .A(net619),
    .B(_0400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3349_ (.A(_0399_),
    .B(_0401_),
    .Y(_0065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3350_ (.B1(net618),
    .VDD(VPWR),
    .Y(_0402_),
    .VSS(VGND),
    .A1(_2585_),
    .A2(_0400_));
 sg13g2_a21oi_1 _3351_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2585_),
    .A2(_0400_),
    .Y(_0066_),
    .B1(_0402_));
 sg13g2_nor2_1 _3352_ (.A(_2584_),
    .B(_0402_),
    .Y(_0067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3353_ (.A(\mydesign.out[0] ),
    .B(\mydesign.out[1] ),
    .X(_0403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3354_ (.S0(net513),
    .A0(\mydesign.accum[96] ),
    .A1(\mydesign.accum[64] ),
    .A2(\mydesign.accum[32] ),
    .A3(\mydesign.accum[0] ),
    .S1(net506),
    .X(_0404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3355_ (.A(net834),
    .B_N(net755),
    .Y(_0405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3356_ (.S0(net515),
    .A0(\mydesign.accum[112] ),
    .A1(\mydesign.accum[80] ),
    .A2(\mydesign.accum[48] ),
    .A3(\mydesign.accum[16] ),
    .S1(net509),
    .X(_0406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3357_ (.A(net755),
    .B(net834),
    .Y(_0407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3358_ (.S0(net511),
    .A0(\mydesign.accum[120] ),
    .A1(\mydesign.accum[88] ),
    .A2(\mydesign.accum[56] ),
    .A3(\mydesign.accum[24] ),
    .S1(net505),
    .X(_0408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3359_ (.A0(\mydesign.accum[104] ),
    .A1(\mydesign.accum[72] ),
    .S(net514),
    .X(_0409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3360_ (.A(net514),
    .B_N(\mydesign.accum[40] ),
    .Y(_0410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3361_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[8] ),
    .A2(net514),
    .Y(_0411_),
    .B1(_0410_));
 sg13g2_nor2b_2 _3362_ (.A(net755),
    .B_N(net834),
    .Y(_0412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3363_ (.B1(_0412_),
    .VDD(VPWR),
    .Y(_0413_),
    .VSS(VGND),
    .A1(net507),
    .A2(_0409_));
 sg13g2_a21oi_1 _3364_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net507),
    .A2(_0411_),
    .Y(_0414_),
    .B1(_0413_));
 sg13g2_a21oi_1 _3365_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net456),
    .A2(_0408_),
    .Y(_0415_),
    .B1(_2698_));
 sg13g2_a221oi_1 _3366_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0406_),
    .C1(_0414_),
    .B1(_0405_),
    .A1(net458),
    .Y(_0416_),
    .A2(_0404_));
 sg13g2_o21ai_1 _3367_ (.B1(net623),
    .VDD(VPWR),
    .Y(_0417_),
    .VSS(VGND),
    .A1(net1081),
    .A2(net430));
 sg13g2_a21oi_1 _3368_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0415_),
    .A2(_0416_),
    .Y(_0068_),
    .B1(_0417_));
 sg13g2_mux4_1 _3369_ (.S0(net513),
    .A0(\mydesign.accum[97] ),
    .A1(\mydesign.accum[65] ),
    .A2(\mydesign.accum[33] ),
    .A3(\mydesign.accum[1] ),
    .S1(net506),
    .X(_0418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3370_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net458),
    .A2(_0418_),
    .Y(_0419_),
    .B1(_2698_));
 sg13g2_mux4_1 _3371_ (.S0(net515),
    .A0(\mydesign.accum[113] ),
    .A1(\mydesign.accum[81] ),
    .A2(\mydesign.accum[49] ),
    .A3(\mydesign.accum[17] ),
    .S1(net508),
    .X(_0420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3372_ (.S0(net511),
    .A0(\mydesign.accum[121] ),
    .A1(\mydesign.accum[89] ),
    .A2(\mydesign.accum[57] ),
    .A3(\mydesign.accum[25] ),
    .S1(net505),
    .X(_0421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3373_ (.A0(\mydesign.accum[105] ),
    .A1(\mydesign.accum[73] ),
    .S(net514),
    .X(_0422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3374_ (.A(net514),
    .B_N(\mydesign.accum[41] ),
    .Y(_0423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3375_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[9] ),
    .A2(net514),
    .Y(_0424_),
    .B1(_0423_));
 sg13g2_o21ai_1 _3376_ (.B1(_0412_),
    .VDD(VPWR),
    .Y(_0425_),
    .VSS(VGND),
    .A1(net507),
    .A2(_0422_));
 sg13g2_a21oi_1 _3377_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net506),
    .A2(_0424_),
    .Y(_0426_),
    .B1(_0425_));
 sg13g2_a221oi_1 _3378_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net456),
    .C1(_0426_),
    .B1(_0421_),
    .A1(_0405_),
    .Y(_0427_),
    .A2(_0420_));
 sg13g2_o21ai_1 _3379_ (.B1(net622),
    .VDD(VPWR),
    .Y(_0428_),
    .VSS(VGND),
    .A1(net1069),
    .A2(net431));
 sg13g2_a21oi_1 _3380_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0419_),
    .A2(_0427_),
    .Y(_0069_),
    .B1(_0428_));
 sg13g2_mux4_1 _3381_ (.S0(net513),
    .A0(\mydesign.accum[106] ),
    .A1(\mydesign.accum[74] ),
    .A2(\mydesign.accum[42] ),
    .A3(\mydesign.accum[10] ),
    .S1(net506),
    .X(_0429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3382_ (.S0(net511),
    .A0(\mydesign.accum[122] ),
    .A1(\mydesign.accum[90] ),
    .A2(\mydesign.accum[58] ),
    .A3(\mydesign.accum[26] ),
    .S1(net505),
    .X(_0430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3383_ (.S0(net515),
    .A0(\mydesign.accum[114] ),
    .A1(\mydesign.accum[82] ),
    .A2(\mydesign.accum[50] ),
    .A3(\mydesign.accum[18] ),
    .S1(net509),
    .X(_0431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3384_ (.A0(\mydesign.accum[98] ),
    .A1(\mydesign.accum[66] ),
    .S(net512),
    .X(_0432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3385_ (.A(net517),
    .B_N(\mydesign.accum[34] ),
    .Y(_0433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3386_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0433_),
    .Y(_0434_),
    .A2(net514),
    .A1(\mydesign.accum[2] ));
 sg13g2_o21ai_1 _3387_ (.B1(net457),
    .VDD(VPWR),
    .Y(_0435_),
    .VSS(VGND),
    .A1(net504),
    .A2(_0432_));
 sg13g2_a21oi_1 _3388_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net504),
    .A2(_0434_),
    .Y(_0436_),
    .B1(_0435_));
 sg13g2_a21oi_1 _3389_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0405_),
    .A2(_0431_),
    .Y(_0437_),
    .B1(_2698_));
 sg13g2_a221oi_1 _3390_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net456),
    .C1(_0436_),
    .B1(_0430_),
    .A1(_0412_),
    .Y(_0438_),
    .A2(_0429_));
 sg13g2_o21ai_1 _3391_ (.B1(net622),
    .VDD(VPWR),
    .Y(_0439_),
    .VSS(VGND),
    .A1(net1087),
    .A2(net430));
 sg13g2_a21oi_1 _3392_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0437_),
    .A2(_0438_),
    .Y(_0070_),
    .B1(_0439_));
 sg13g2_mux4_1 _3393_ (.S0(net515),
    .A0(\mydesign.accum[115] ),
    .A1(\mydesign.accum[83] ),
    .A2(\mydesign.accum[51] ),
    .A3(\mydesign.accum[19] ),
    .S1(net508),
    .X(_0440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3394_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0405_),
    .A2(_0440_),
    .Y(_0441_),
    .B1(_2698_));
 sg13g2_mux4_1 _3395_ (.S0(net511),
    .A0(\mydesign.accum[123] ),
    .A1(\mydesign.accum[91] ),
    .A2(\mydesign.accum[59] ),
    .A3(\mydesign.accum[27] ),
    .S1(net504),
    .X(_0442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3396_ (.S0(net513),
    .A0(\mydesign.accum[107] ),
    .A1(\mydesign.accum[75] ),
    .A2(\mydesign.accum[43] ),
    .A3(\mydesign.accum[11] ),
    .S1(net506),
    .X(_0443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3397_ (.A0(\mydesign.accum[99] ),
    .A1(\mydesign.accum[67] ),
    .S(net512),
    .X(_0444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3398_ (.A(net517),
    .B_N(\mydesign.accum[35] ),
    .Y(_0445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3399_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0445_),
    .Y(_0446_),
    .A2(net517),
    .A1(\mydesign.accum[3] ));
 sg13g2_o21ai_1 _3400_ (.B1(net458),
    .VDD(VPWR),
    .Y(_0447_),
    .VSS(VGND),
    .A1(net504),
    .A2(_0444_));
 sg13g2_a21oi_1 _3401_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net504),
    .A2(_0446_),
    .Y(_0448_),
    .B1(_0447_));
 sg13g2_a221oi_1 _3402_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0412_),
    .C1(_0448_),
    .B1(_0443_),
    .A1(net456),
    .Y(_0449_),
    .A2(_0442_));
 sg13g2_o21ai_1 _3403_ (.B1(net627),
    .VDD(VPWR),
    .Y(_0450_),
    .VSS(VGND),
    .A1(net1078),
    .A2(net430));
 sg13g2_a21oi_1 _3404_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0441_),
    .A2(_0449_),
    .Y(_0071_),
    .B1(_0450_));
 sg13g2_mux4_1 _3405_ (.S0(net513),
    .A0(\mydesign.accum[108] ),
    .A1(\mydesign.accum[76] ),
    .A2(\mydesign.accum[44] ),
    .A3(\mydesign.accum[12] ),
    .S1(net508),
    .X(_0451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3406_ (.S0(net518),
    .A0(\mydesign.accum[124] ),
    .A1(\mydesign.accum[92] ),
    .A2(\mydesign.accum[60] ),
    .A3(\mydesign.accum[28] ),
    .S1(net505),
    .X(_0452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3407_ (.S0(net515),
    .A0(\mydesign.accum[116] ),
    .A1(\mydesign.accum[84] ),
    .A2(\mydesign.accum[52] ),
    .A3(\mydesign.accum[20] ),
    .S1(net508),
    .X(_0453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3408_ (.S0(net512),
    .A0(\mydesign.accum[100] ),
    .A1(\mydesign.accum[68] ),
    .A2(\mydesign.accum[36] ),
    .A3(\mydesign.accum[4] ),
    .S1(net507),
    .X(_0454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3409_ (.Y(_0455_),
    .B1(_0454_),
    .B2(net457),
    .A2(_0452_),
    .A1(net456),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3410_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0405_),
    .C1(_2698_),
    .B1(_0453_),
    .A1(_0412_),
    .Y(_0456_),
    .A2(_0451_));
 sg13g2_o21ai_1 _3411_ (.B1(net622),
    .VDD(VPWR),
    .Y(_0457_),
    .VSS(VGND),
    .A1(net1075),
    .A2(net430));
 sg13g2_a21oi_1 _3412_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0455_),
    .A2(_0456_),
    .Y(_0072_),
    .B1(_0457_));
 sg13g2_mux2_1 _3413_ (.A0(\mydesign.accum[125] ),
    .A1(\mydesign.accum[93] ),
    .S(net511),
    .X(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3414_ (.B1(net505),
    .VDD(VPWR),
    .Y(_0459_),
    .VSS(VGND),
    .A1(_2548_),
    .A2(net511));
 sg13g2_a21oi_1 _3415_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net890),
    .A2(net512),
    .Y(_0460_),
    .B1(_0459_));
 sg13g2_o21ai_1 _3416_ (.B1(_0407_),
    .VDD(VPWR),
    .Y(_0461_),
    .VSS(VGND),
    .A1(net504),
    .A2(_0458_));
 sg13g2_o21ai_1 _3417_ (.B1(net430),
    .VDD(VPWR),
    .Y(_0462_),
    .VSS(VGND),
    .A1(_0460_),
    .A2(_0461_));
 sg13g2_mux4_1 _3418_ (.S0(net516),
    .A0(\mydesign.accum[117] ),
    .A1(\mydesign.accum[85] ),
    .A2(\mydesign.accum[53] ),
    .A3(\mydesign.accum[21] ),
    .S1(net508),
    .X(_0463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3419_ (.S0(net515),
    .A0(\mydesign.accum[109] ),
    .A1(\mydesign.accum[77] ),
    .A2(\mydesign.accum[45] ),
    .A3(\mydesign.accum[13] ),
    .S1(net508),
    .X(_0464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3420_ (.S0(net513),
    .A0(\mydesign.accum[101] ),
    .A1(\mydesign.accum[69] ),
    .A2(\mydesign.accum[37] ),
    .A3(\mydesign.accum[5] ),
    .S1(net506),
    .X(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3421_ (.Y(_0466_),
    .B1(_0464_),
    .B2(_0412_),
    .A2(_0463_),
    .A1(_0405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3422_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net457),
    .A2(_0465_),
    .Y(_0467_),
    .B1(_0462_));
 sg13g2_o21ai_1 _3423_ (.B1(net622),
    .VDD(VPWR),
    .Y(_0468_),
    .VSS(VGND),
    .A1(net1080),
    .A2(net431));
 sg13g2_a21oi_1 _3424_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0466_),
    .A2(_0467_),
    .Y(_0073_),
    .B1(_0468_));
 sg13g2_mux4_1 _3425_ (.S0(net511),
    .A0(\mydesign.accum[126] ),
    .A1(\mydesign.accum[94] ),
    .A2(\mydesign.accum[62] ),
    .A3(\mydesign.accum[30] ),
    .S1(net505),
    .X(_0469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3426_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net456),
    .A2(_0469_),
    .Y(_0470_),
    .B1(_2698_));
 sg13g2_mux4_1 _3427_ (.S0(net515),
    .A0(\mydesign.accum[110] ),
    .A1(\mydesign.accum[78] ),
    .A2(\mydesign.accum[46] ),
    .A3(\mydesign.accum[14] ),
    .S1(net508),
    .X(_0471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3428_ (.S0(net513),
    .A0(\mydesign.accum[102] ),
    .A1(\mydesign.accum[70] ),
    .A2(\mydesign.accum[38] ),
    .A3(\mydesign.accum[6] ),
    .S1(net506),
    .X(_0472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3429_ (.A0(\mydesign.accum[118] ),
    .A1(\mydesign.accum[86] ),
    .S(net512),
    .X(_0473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3430_ (.A(net516),
    .B_N(\mydesign.accum[54] ),
    .Y(_0474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3431_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[22] ),
    .A2(net516),
    .Y(_0475_),
    .B1(_0474_));
 sg13g2_o21ai_1 _3432_ (.B1(_0405_),
    .VDD(VPWR),
    .Y(_0476_),
    .VSS(VGND),
    .A1(net509),
    .A2(_0473_));
 sg13g2_a21oi_1 _3433_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net509),
    .A2(_0475_),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_a221oi_1 _3434_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net458),
    .C1(_0477_),
    .B1(_0472_),
    .A1(_0412_),
    .Y(_0478_),
    .A2(_0471_));
 sg13g2_o21ai_1 _3435_ (.B1(net622),
    .VDD(VPWR),
    .Y(_0479_),
    .VSS(VGND),
    .A1(net1072),
    .A2(net430));
 sg13g2_a21oi_1 _3436_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0470_),
    .A2(_0478_),
    .Y(_0074_),
    .B1(_0479_));
 sg13g2_mux4_1 _3437_ (.S0(net515),
    .A0(\mydesign.accum[111] ),
    .A1(\mydesign.accum[79] ),
    .A2(\mydesign.accum[47] ),
    .A3(\mydesign.accum[15] ),
    .S1(net508),
    .X(_0480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3438_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0412_),
    .A2(_0480_),
    .Y(_0481_),
    .B1(_2698_));
 sg13g2_mux4_1 _3439_ (.S0(net513),
    .A0(\mydesign.accum[103] ),
    .A1(\mydesign.accum[71] ),
    .A2(\mydesign.accum[39] ),
    .A3(\mydesign.accum[7] ),
    .S1(net506),
    .X(_0482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3440_ (.S0(net511),
    .A0(\mydesign.accum[127] ),
    .A1(\mydesign.accum[95] ),
    .A2(\mydesign.accum[63] ),
    .A3(\mydesign.accum[31] ),
    .S1(net505),
    .X(_0483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3441_ (.A0(\mydesign.accum[119] ),
    .A1(\mydesign.accum[87] ),
    .S(net516),
    .X(_0484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3442_ (.A(net516),
    .B_N(\mydesign.accum[55] ),
    .Y(_0485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3443_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[23] ),
    .A2(net516),
    .Y(_0486_),
    .B1(_0485_));
 sg13g2_o21ai_1 _3444_ (.B1(_0405_),
    .VDD(VPWR),
    .Y(_0487_),
    .VSS(VGND),
    .A1(net509),
    .A2(_0484_));
 sg13g2_a21oi_1 _3445_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net509),
    .A2(_0486_),
    .Y(_0488_),
    .B1(_0487_));
 sg13g2_a221oi_1 _3446_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net456),
    .C1(_0488_),
    .B1(_0483_),
    .A1(net457),
    .Y(_0489_),
    .A2(_0482_));
 sg13g2_o21ai_1 _3447_ (.B1(net622),
    .VDD(VPWR),
    .Y(_0490_),
    .VSS(VGND),
    .A1(net1084),
    .A2(net430));
 sg13g2_a21oi_1 _3448_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0481_),
    .A2(_0489_),
    .Y(_0075_),
    .B1(_0490_));
 sg13g2_nor2_1 _3449_ (.A(_2639_),
    .B(_2683_),
    .Y(_0491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3450_ (.Y(_0492_),
    .A(net606),
    .B(_0491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3451_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net607),
    .Y(_0493_),
    .A2(_0491_),
    .A1(net606));
 sg13g2_nand2_1 _3452_ (.Y(_0494_),
    .A(net414),
    .B(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3453_ (.B1(_0494_),
    .VDD(VPWR),
    .Y(_0076_),
    .VSS(VGND),
    .A1(net604),
    .A2(_0492_));
 sg13g2_nand2_1 _3454_ (.Y(_0495_),
    .A(net425),
    .B(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3455_ (.B1(_0495_),
    .VDD(VPWR),
    .Y(_0077_),
    .VSS(VGND),
    .A1(net602),
    .A2(_0492_));
 sg13g2_nand2_1 _3456_ (.Y(_0496_),
    .A(net418),
    .B(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3457_ (.B1(_0496_),
    .VDD(VPWR),
    .Y(_0078_),
    .VSS(VGND),
    .A1(net599),
    .A2(_0492_));
 sg13g2_nand2_1 _3458_ (.Y(_0497_),
    .A(net652),
    .B(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3459_ (.B1(_0497_),
    .VDD(VPWR),
    .Y(_0079_),
    .VSS(VGND),
    .A1(net597),
    .A2(_0492_));
 sg13g2_mux4_1 _3460_ (.S0(net554),
    .A0(\mydesign.inputs[0][24] ),
    .A1(\mydesign.inputs[0][20] ),
    .A2(\mydesign.inputs[0][16] ),
    .A3(\mydesign.inputs[0][12] ),
    .S1(net544),
    .X(_0498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3461_ (.A(net542),
    .B(net484),
    .Y(_0499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3462_ (.Y(_0500_),
    .B1(net455),
    .B2(_0499_),
    .A2(net484),
    .A1(net540),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3463_ (.A(net609),
    .B(_0500_),
    .Y(_0080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3464_ (.S0(net554),
    .A0(\mydesign.inputs[0][25] ),
    .A1(\mydesign.inputs[0][21] ),
    .A2(\mydesign.inputs[0][17] ),
    .A3(\mydesign.inputs[0][13] ),
    .S1(net544),
    .X(_0501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3465_ (.Y(_0502_),
    .B1(_0499_),
    .B2(_0501_),
    .A2(net484),
    .A1(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3466_ (.A(net609),
    .B(_0502_),
    .Y(_0081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3467_ (.A(net554),
    .B_N(\mydesign.inputs[0][26] ),
    .Y(_0503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3468_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net554),
    .A2(\mydesign.inputs[0][22] ),
    .Y(_0504_),
    .B1(_0503_));
 sg13g2_a22oi_1 _3469_ (.Y(_0505_),
    .B1(_0394_),
    .B2(\mydesign.inputs[0][14] ),
    .A2(net495),
    .A1(\mydesign.inputs[0][18] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3470_ (.B1(_0505_),
    .VDD(VPWR),
    .Y(_0506_),
    .VSS(VGND),
    .A1(net544),
    .A2(_0504_));
 sg13g2_a21oi_1 _3471_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2586_),
    .A2(_0506_),
    .Y(_0507_),
    .B1(net484));
 sg13g2_o21ai_1 _3472_ (.B1(net627),
    .VDD(VPWR),
    .Y(_0508_),
    .VSS(VGND),
    .A1(net1086),
    .A2(net436));
 sg13g2_nor2_1 _3473_ (.A(_0507_),
    .B(_0508_),
    .Y(_0082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3474_ (.A(net554),
    .B_N(\mydesign.inputs[0][27] ),
    .Y(_0509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3475_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net554),
    .A2(\mydesign.inputs[0][23] ),
    .Y(_0510_),
    .B1(_0509_));
 sg13g2_a22oi_1 _3476_ (.Y(_0511_),
    .B1(_0394_),
    .B2(\mydesign.inputs[0][15] ),
    .A2(net495),
    .A1(\mydesign.inputs[0][19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3477_ (.B1(_0511_),
    .VDD(VPWR),
    .Y(_0512_),
    .VSS(VGND),
    .A1(net544),
    .A2(_0510_));
 sg13g2_a22oi_1 _3478_ (.Y(_0513_),
    .B1(_0499_),
    .B2(_0512_),
    .A2(net484),
    .A1(net1059),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3479_ (.A(net609),
    .B(_0513_),
    .Y(_0083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3480_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net498),
    .A2(_2592_),
    .Y(_0514_),
    .B1(net546));
 sg13g2_o21ai_1 _3481_ (.B1(_0514_),
    .VDD(VPWR),
    .Y(_0515_),
    .VSS(VGND),
    .A1(net498),
    .A2(\mydesign.weights[0][20] ));
 sg13g2_a22oi_1 _3482_ (.Y(_0516_),
    .B1(_0394_),
    .B2(\mydesign.weights[0][12] ),
    .A2(net496),
    .A1(\mydesign.weights[0][16] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3483_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net543),
    .Y(_0517_),
    .A2(_0516_),
    .A1(_0515_));
 sg13g2_o21ai_1 _3484_ (.B1(net621),
    .VDD(VPWR),
    .Y(_0518_),
    .VSS(VGND),
    .A1(net485),
    .A2(_0517_));
 sg13g2_a21oi_1 _3485_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2578_),
    .A2(net484),
    .Y(_0084_),
    .B1(_0518_));
 sg13g2_mux4_1 _3486_ (.S0(net553),
    .A0(\mydesign.weights[0][25] ),
    .A1(\mydesign.weights[0][21] ),
    .A2(\mydesign.weights[0][17] ),
    .A3(\mydesign.weights[0][13] ),
    .S1(net546),
    .X(_0519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3487_ (.A(_2586_),
    .B(_0519_),
    .X(_0520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3488_ (.B1(net621),
    .VDD(VPWR),
    .Y(_0521_),
    .VSS(VGND),
    .A1(net485),
    .A2(_0520_));
 sg13g2_a21oi_1 _3489_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2577_),
    .A2(net484),
    .Y(_0085_),
    .B1(_0521_));
 sg13g2_mux4_1 _3490_ (.S0(net553),
    .A0(\mydesign.weights[0][26] ),
    .A1(\mydesign.weights[0][22] ),
    .A2(\mydesign.weights[0][18] ),
    .A3(\mydesign.weights[0][14] ),
    .S1(net546),
    .X(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3491_ (.A(_2586_),
    .B(_0522_),
    .X(_0523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3492_ (.B1(net624),
    .VDD(VPWR),
    .Y(_0524_),
    .VSS(VGND),
    .A1(net485),
    .A2(_0523_));
 sg13g2_a21oi_1 _3493_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2576_),
    .A2(net485),
    .Y(_0086_),
    .B1(_0524_));
 sg13g2_mux4_1 _3494_ (.S0(net556),
    .A0(\mydesign.weights[0][27] ),
    .A1(\mydesign.weights[0][23] ),
    .A2(\mydesign.weights[0][19] ),
    .A3(\mydesign.weights[0][15] ),
    .S1(net545),
    .X(_0525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3495_ (.A(_2586_),
    .B(_0525_),
    .X(_0526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3496_ (.B1(net624),
    .VDD(VPWR),
    .Y(_0527_),
    .VSS(VGND),
    .A1(net484),
    .A2(_0526_));
 sg13g2_a21oi_1 _3497_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2575_),
    .A2(net485),
    .Y(_0087_),
    .B1(_0527_));
 sg13g2_and3_1 _3498_ (.X(_0528_),
    .A(net558),
    .B(net455),
    .C(_0517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3499_ (.B1(net467),
    .VDD(VPWR),
    .Y(_0529_),
    .VSS(VGND),
    .A1(net721),
    .A2(_0528_));
 sg13g2_a21oi_1 _3500_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net721),
    .A2(_0528_),
    .Y(_0088_),
    .B1(_0529_));
 sg13g2_nand3_1 _3501_ (.B(net455),
    .C(_0520_),
    .A(\mydesign.accum[121] ),
    .Y(_0530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3502_ (.A2(_0520_),
    .A1(net455),
    .B1(\mydesign.accum[121] ),
    .X(_0531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3503_ (.Y(_0532_),
    .A(_0530_),
    .B(_0531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3504_ (.Y(_0533_),
    .A(_0501_),
    .B(_0517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3505_ (.A(_0532_),
    .B(_0533_),
    .Y(_0534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3506_ (.B(_0533_),
    .A(_0532_),
    .X(_0535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3507_ (.B(net455),
    .C(_0517_),
    .A(net721),
    .Y(_0536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3508_ (.B(net455),
    .C(_0517_),
    .A(net721),
    .Y(_0537_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0535_));
 sg13g2_xor2_1 _3509_ (.B(_0536_),
    .A(_0535_),
    .X(_0538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3510_ (.B1(net467),
    .VDD(VPWR),
    .Y(_0539_),
    .VSS(VGND),
    .A1(net558),
    .A2(net937));
 sg13g2_a21oi_1 _3511_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net558),
    .A2(_0538_),
    .Y(_0089_),
    .B1(_0539_));
 sg13g2_nand2_1 _3512_ (.Y(_0540_),
    .A(_0506_),
    .B(_0517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3513_ (.B(net455),
    .C(_0523_),
    .A(\mydesign.accum[122] ),
    .Y(_0541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3514_ (.A2(_0523_),
    .A1(_0498_),
    .B1(\mydesign.accum[122] ),
    .X(_0542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3515_ (.Y(_0543_),
    .A(_0541_),
    .B(_0542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3516_ (.Y(_0544_),
    .A(_0501_),
    .B(_0520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3517_ (.A(_0543_),
    .B(_0544_),
    .Y(_0545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3518_ (.B(_0544_),
    .A(_0543_),
    .X(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3519_ (.Y(_0547_),
    .B(_0546_),
    .A_N(_0530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3520_ (.Y(_0548_),
    .A(_0530_),
    .B(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3521_ (.Y(_0549_),
    .B(_0548_),
    .A_N(_0540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3522_ (.Y(_0550_),
    .A(_0540_),
    .B(_0548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3523_ (.Y(_0551_),
    .A(_0534_),
    .B(_0550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3524_ (.Y(_0552_),
    .A(_0534_),
    .B(_0550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3525_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0553_),
    .B(_0552_),
    .A(_0537_));
 sg13g2_xnor2_1 _3526_ (.Y(_0554_),
    .A(_0537_),
    .B(_0552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3527_ (.B1(net467),
    .VDD(VPWR),
    .Y(_0555_),
    .VSS(VGND),
    .A1(net558),
    .A2(net958));
 sg13g2_a21oi_1 _3528_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net558),
    .A2(_0554_),
    .Y(_0090_),
    .B1(_0555_));
 sg13g2_nand2_1 _3529_ (.Y(_0556_),
    .A(_0547_),
    .B(_0549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3530_ (.Y(_0557_),
    .A(_0512_),
    .B(_0517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3531_ (.Y(_0558_),
    .A(_0506_),
    .B(_0520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3532_ (.Y(_0559_),
    .A(_0501_),
    .B(_0523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3533_ (.B(net455),
    .C(_0525_),
    .A(_2586_),
    .Y(_0560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3534_ (.B(_0498_),
    .C(_0526_),
    .A(\mydesign.accum[123] ),
    .Y(_0561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3535_ (.B(_0560_),
    .A(\mydesign.accum[123] ),
    .X(_0562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3536_ (.B(_0562_),
    .A(_0559_),
    .X(_0563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3537_ (.Y(_0564_),
    .B(_0563_),
    .A_N(_0541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3538_ (.Y(_0565_),
    .A(_0541_),
    .B(_0563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3539_ (.Y(_0566_),
    .B(_0565_),
    .A_N(_0558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3540_ (.Y(_0567_),
    .A(_0558_),
    .B(_0565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3541_ (.Y(_0568_),
    .A(_0545_),
    .B(_0567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3542_ (.A(_0545_),
    .B(_0567_),
    .Y(_0569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3543_ (.B(_0567_),
    .A(_0545_),
    .X(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3544_ (.Y(_0571_),
    .A(_0557_),
    .B(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3545_ (.Y(_0572_),
    .A(_0556_),
    .B(_0571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3546_ (.Y(_0573_),
    .A(_0556_),
    .B(_0571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3547_ (.B(_0553_),
    .C(_0573_),
    .A(_0551_),
    .Y(_0574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3548_ (.A2(_0553_),
    .A1(_0551_),
    .B1(_0573_),
    .X(_0575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3549_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0574_),
    .A2(_0575_),
    .Y(_0576_),
    .B1(net499));
 sg13g2_o21ai_1 _3550_ (.B1(net468),
    .VDD(VPWR),
    .Y(_0577_),
    .VSS(VGND),
    .A1(net559),
    .A2(net1061));
 sg13g2_nor2_1 _3551_ (.A(_0576_),
    .B(_0577_),
    .Y(_0091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3552_ (.Y(_0578_),
    .A(_0564_),
    .B(_0566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3553_ (.Y(_0579_),
    .A(_0512_),
    .B(_0520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3554_ (.B1(_0561_),
    .VDD(VPWR),
    .Y(_0580_),
    .VSS(VGND),
    .A1(_0559_),
    .A2(_0562_));
 sg13g2_nand2_1 _3555_ (.Y(_0581_),
    .A(_0506_),
    .B(_0523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3556_ (.B(_0501_),
    .C(_0526_),
    .A(\mydesign.accum[124] ),
    .Y(_0582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3557_ (.A2(_0526_),
    .A1(_0501_),
    .B1(\mydesign.accum[124] ),
    .X(_0583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3558_ (.Y(_0584_),
    .A(_0582_),
    .B(_0583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3559_ (.B(_0584_),
    .A(_0581_),
    .X(_0585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3560_ (.Y(_0586_),
    .A(_0580_),
    .B(_0585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3561_ (.Y(_0587_),
    .A(_0580_),
    .B(_0585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3562_ (.B(_0587_),
    .A(_0579_),
    .X(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3563_ (.Y(_0589_),
    .A(_0578_),
    .B(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3564_ (.Y(_0590_),
    .A(_0578_),
    .B(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3565_ (.B1(_0568_),
    .VDD(VPWR),
    .Y(_0591_),
    .VSS(VGND),
    .A1(_0557_),
    .A2(_0569_));
 sg13g2_nand2b_1 _3566_ (.Y(_0592_),
    .B(_0591_),
    .A_N(_0590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3567_ (.B(_0591_),
    .A(_0590_),
    .X(_0593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3568_ (.B(_0575_),
    .C(_0593_),
    .A(_0572_),
    .Y(_0594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3569_ (.A2(_0575_),
    .A1(_0572_),
    .B1(_0593_),
    .X(_0595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3570_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0594_),
    .A2(_0595_),
    .Y(_0596_),
    .B1(net500));
 sg13g2_o21ai_1 _3571_ (.B1(net468),
    .VDD(VPWR),
    .Y(_0597_),
    .VSS(VGND),
    .A1(net559),
    .A2(net1079));
 sg13g2_nor2_1 _3572_ (.A(_0596_),
    .B(_0597_),
    .Y(_0092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3573_ (.Y(_0598_),
    .A(_0592_),
    .B(_0595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3574_ (.B1(_0586_),
    .VDD(VPWR),
    .Y(_0599_),
    .VSS(VGND),
    .A1(_0579_),
    .A2(_0587_));
 sg13g2_nand2_1 _3575_ (.Y(_0600_),
    .A(_0512_),
    .B(_0523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3576_ (.A(_0506_),
    .B(_0526_),
    .X(_0601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3577_ (.Y(_0602_),
    .A(\mydesign.accum[125] ),
    .B(_0601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3578_ (.A(_0600_),
    .B(_0602_),
    .Y(_0603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3579_ (.B(_0602_),
    .A(_0600_),
    .X(_0604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3580_ (.B1(_0582_),
    .VDD(VPWR),
    .Y(_0605_),
    .VSS(VGND),
    .A1(_0581_),
    .A2(_0584_));
 sg13g2_nand2_1 _3581_ (.Y(_0606_),
    .A(_0604_),
    .B(_0605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3582_ (.B(_0605_),
    .A(_0604_),
    .X(_0607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3583_ (.Y(_0608_),
    .A(_0599_),
    .B(_0607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3584_ (.Y(_0609_),
    .A(_0599_),
    .B(_0607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3585_ (.A(_0589_),
    .B(_0609_),
    .Y(_0610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3586_ (.Y(_0611_),
    .A(_0589_),
    .B(_0609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3587_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0592_),
    .A2(_0595_),
    .Y(_0612_),
    .B1(_0611_));
 sg13g2_xor2_1 _3588_ (.B(_0611_),
    .A(_0598_),
    .X(_0613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3589_ (.B1(net468),
    .VDD(VPWR),
    .Y(_0614_),
    .VSS(VGND),
    .A1(net558),
    .A2(net1060));
 sg13g2_a21oi_1 _3590_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net558),
    .A2(_0613_),
    .Y(_0093_),
    .B1(_0614_));
 sg13g2_a21oi_1 _3591_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[125] ),
    .A2(_0601_),
    .Y(_0615_),
    .B1(_0603_));
 sg13g2_nand3_1 _3592_ (.B(_0512_),
    .C(_0526_),
    .A(\mydesign.accum[126] ),
    .Y(_0616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3593_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0512_),
    .A2(_0526_),
    .Y(_0617_),
    .B1(\mydesign.accum[126] ));
 sg13g2_a21o_1 _3594_ (.A2(_0526_),
    .A1(_0512_),
    .B1(\mydesign.accum[126] ),
    .X(_0618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3595_ (.Y(_0619_),
    .A(_0616_),
    .B(_0618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3596_ (.Y(_0620_),
    .A(_0615_),
    .B(_0619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3597_ (.A(_0606_),
    .B(_0620_),
    .Y(_0621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3598_ (.B(_0620_),
    .A(_0606_),
    .X(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3599_ (.Y(_0623_),
    .B(_0622_),
    .A_N(_0608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3600_ (.Y(_0624_),
    .A(_0608_),
    .B(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3601_ (.A(_0610_),
    .B(_0612_),
    .C(_0624_),
    .X(_0625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3602_ (.B1(_0624_),
    .VDD(VPWR),
    .Y(_0626_),
    .VSS(VGND),
    .A1(_0610_),
    .A2(_0612_));
 sg13g2_a21oi_1 _3603_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0625_),
    .A2(_0626_),
    .Y(_0627_),
    .B1(net500));
 sg13g2_o21ai_1 _3604_ (.B1(net468),
    .VDD(VPWR),
    .Y(_0628_),
    .VSS(VGND),
    .A1(net558),
    .A2(net1062));
 sg13g2_nor2_1 _3605_ (.A(_0627_),
    .B(_0628_),
    .Y(_0094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3606_ (.Y(_0629_),
    .A(_0623_),
    .B(_0626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3607_ (.B1(_0616_),
    .VDD(VPWR),
    .Y(_0630_),
    .VSS(VGND),
    .A1(_0615_),
    .A2(_0617_));
 sg13g2_xnor2_1 _3608_ (.Y(_0631_),
    .A(net1004),
    .B(_0630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3609_ (.Y(_0632_),
    .A(_0621_),
    .B(_0631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3610_ (.Y(_0633_),
    .A(_0629_),
    .B(_0632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3611_ (.B1(net468),
    .VDD(VPWR),
    .Y(_0634_),
    .VSS(VGND),
    .A1(net559),
    .A2(net1004));
 sg13g2_a21oi_1 _3612_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net559),
    .A2(_0633_),
    .Y(_0095_),
    .B1(_0634_));
 sg13g2_o21ai_1 _3613_ (.B1(net626),
    .VDD(VPWR),
    .Y(_0635_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[60] ),
    .A2(net487));
 sg13g2_a21oi_1 _3614_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2583_),
    .A2(net486),
    .Y(_0096_),
    .B1(_0635_));
 sg13g2_o21ai_1 _3615_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0636_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[61] ),
    .A2(net487));
 sg13g2_a21oi_1 _3616_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2582_),
    .A2(net486),
    .Y(_0097_),
    .B1(_0636_));
 sg13g2_o21ai_1 _3617_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0637_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[62] ),
    .A2(net487));
 sg13g2_a21oi_1 _3618_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2581_),
    .A2(net490),
    .Y(_0098_),
    .B1(_0637_));
 sg13g2_o21ai_1 _3619_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0638_),
    .VSS(VGND),
    .A1(net1059),
    .A2(net487));
 sg13g2_a21oi_1 _3620_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2580_),
    .A2(net490),
    .Y(_0099_),
    .B1(_0638_));
 sg13g2_nor2_2 _3621_ (.A(net556),
    .B(_0397_),
    .Y(_0639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3622_ (.Y(_0640_),
    .A(\mydesign.weights[1][16] ),
    .B(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3623_ (.Y(_0641_),
    .B1(_0394_),
    .B2(\mydesign.weights[1][12] ),
    .A2(net461),
    .A1(\mydesign.weights[1][20] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3624_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0640_),
    .A2(_0641_),
    .Y(_0642_),
    .B1(net542));
 sg13g2_a21o_2 _3625_ (.A2(_0639_),
    .A1(net802),
    .B1(_0642_),
    .X(_0643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3626_ (.B1(net626),
    .VDD(VPWR),
    .Y(_0644_),
    .VSS(VGND),
    .A1(net487),
    .A2(_0643_));
 sg13g2_a21oi_1 _3627_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2567_),
    .A2(net488),
    .Y(_0100_),
    .B1(_0644_));
 sg13g2_nand2_1 _3628_ (.Y(_0645_),
    .A(\mydesign.weights[1][13] ),
    .B(_0394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3629_ (.Y(_0646_),
    .B1(net461),
    .B2(\mydesign.weights[1][21] ),
    .A2(net495),
    .A1(\mydesign.weights[1][17] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3630_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0645_),
    .A2(_0646_),
    .Y(_0647_),
    .B1(net542));
 sg13g2_a21o_2 _3631_ (.A2(_0639_),
    .A1(net774),
    .B1(_0647_),
    .X(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3632_ (.B1(net631),
    .VDD(VPWR),
    .Y(_0649_),
    .VSS(VGND),
    .A1(net492),
    .A2(_0648_));
 sg13g2_a21oi_1 _3633_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2566_),
    .A2(net492),
    .Y(_0101_),
    .B1(_0649_));
 sg13g2_nand3_1 _3634_ (.B(\mydesign.weights[1][10] ),
    .C(net460),
    .A(net498),
    .Y(_0650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3635_ (.X(_0651_),
    .A(net545),
    .B(net556),
    .C(\mydesign.weights[1][14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3636_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\mydesign.weights[1][22] ),
    .C1(_0651_),
    .B1(net461),
    .A1(\mydesign.weights[1][18] ),
    .Y(_0652_),
    .A2(net495));
 sg13g2_o21ai_1 _3637_ (.B1(_0650_),
    .VDD(VPWR),
    .Y(_0653_),
    .VSS(VGND),
    .A1(net542),
    .A2(_0652_));
 sg13g2_o21ai_1 _3638_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0654_),
    .VSS(VGND),
    .A1(net487),
    .A2(_0653_));
 sg13g2_a21oi_1 _3639_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2565_),
    .A2(net492),
    .Y(_0102_),
    .B1(_0654_));
 sg13g2_nand3_1 _3640_ (.B(\mydesign.weights[1][11] ),
    .C(net460),
    .A(net498),
    .Y(_0655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3641_ (.X(_0656_),
    .A(net545),
    .B(net555),
    .C(\mydesign.weights[1][15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3642_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\mydesign.weights[1][23] ),
    .C1(_0656_),
    .B1(net461),
    .A1(\mydesign.weights[1][19] ),
    .Y(_0657_),
    .A2(net495));
 sg13g2_o21ai_1 _3643_ (.B1(_0655_),
    .VDD(VPWR),
    .Y(_0658_),
    .VSS(VGND),
    .A1(net542),
    .A2(_0657_));
 sg13g2_o21ai_1 _3644_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0659_),
    .VSS(VGND),
    .A1(net492),
    .A2(_0658_));
 sg13g2_a21oi_1 _3645_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2564_),
    .A2(net492),
    .Y(_0103_),
    .B1(_0659_));
 sg13g2_and2_1 _3646_ (.A(net540),
    .B(_0643_),
    .X(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3647_ (.Y(_0661_),
    .A(net577),
    .B(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3648_ (.B(_0661_),
    .A(net991),
    .X(_0662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3649_ (.A(net463),
    .B(_0662_),
    .Y(_0104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3650_ (.B(net540),
    .C(_0648_),
    .A(\mydesign.accum[113] ),
    .Y(_0663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3651_ (.VDD(VPWR),
    .Y(_0664_),
    .A(_0663_),
    .VSS(VGND));
 sg13g2_a21o_1 _3652_ (.A2(_0648_),
    .A1(net540),
    .B1(\mydesign.accum[113] ),
    .X(_0665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3653_ (.A(\mydesign.pe_inputs[61] ),
    .B(_0643_),
    .C(_0663_),
    .D(_0665_),
    .X(_0666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3654_ (.Y(_0667_),
    .B1(_0663_),
    .B2(_0665_),
    .A2(_0643_),
    .A1(\mydesign.pe_inputs[61] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3655_ (.A(_0666_),
    .B(_0667_),
    .Y(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3656_ (.B(_0660_),
    .C(_0668_),
    .A(\mydesign.accum[112] ),
    .Y(_0669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3657_ (.A2(_0660_),
    .A1(\mydesign.accum[112] ),
    .B1(_0668_),
    .X(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3658_ (.Y(_0671_),
    .A(_0669_),
    .B(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3659_ (.B1(net480),
    .VDD(VPWR),
    .Y(_0672_),
    .VSS(VGND),
    .A1(net578),
    .A2(net851));
 sg13g2_a21oi_1 _3660_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net578),
    .A2(_0671_),
    .Y(_0105_),
    .B1(_0672_));
 sg13g2_nand2_1 _3661_ (.Y(_0673_),
    .A(\mydesign.pe_inputs[62] ),
    .B(_0643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3662_ (.X(_0674_),
    .A(\mydesign.accum[114] ),
    .B(net540),
    .C(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3663_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net540),
    .A2(_0653_),
    .Y(_0675_),
    .B1(\mydesign.accum[114] ));
 sg13g2_nor2_1 _3664_ (.A(_0674_),
    .B(_0675_),
    .Y(_0676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3665_ (.Y(_0677_),
    .A(\mydesign.pe_inputs[61] ),
    .B(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3666_ (.A(_0674_),
    .B(_0675_),
    .C(_0677_),
    .Y(_0678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3667_ (.Y(_0679_),
    .A(_0676_),
    .B(_0677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3668_ (.Y(_0680_),
    .A(_0663_),
    .B(_0679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3669_ (.A(_0673_),
    .B_N(_0680_),
    .Y(_0681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3670_ (.Y(_0682_),
    .A(_0673_),
    .B(_0680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3671_ (.Y(_0683_),
    .A(_0666_),
    .B(_0682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3672_ (.Y(_0684_),
    .A(_0666_),
    .B(_0682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3673_ (.Y(_0685_),
    .A(_0669_),
    .B(_0684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3674_ (.B1(net470),
    .VDD(VPWR),
    .Y(_0686_),
    .VSS(VGND),
    .A1(net577),
    .A2(net877));
 sg13g2_a21oi_1 _3675_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net577),
    .A2(_0685_),
    .Y(_0106_),
    .B1(_0686_));
 sg13g2_o21ai_1 _3676_ (.B1(_0683_),
    .VDD(VPWR),
    .Y(_0687_),
    .VSS(VGND),
    .A1(_0669_),
    .A2(_0684_));
 sg13g2_a21oi_1 _3677_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0664_),
    .A2(_0679_),
    .Y(_0688_),
    .B1(_0681_));
 sg13g2_and2_1 _3678_ (.A(\mydesign.pe_inputs[63] ),
    .B(_0643_),
    .X(_0689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3679_ (.Y(_0690_),
    .A(\mydesign.pe_inputs[62] ),
    .B(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3680_ (.Y(_0691_),
    .A(\mydesign.pe_inputs[61] ),
    .B(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3681_ (.X(_0692_),
    .A(\mydesign.accum[115] ),
    .B(net540),
    .C(_0658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3682_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net540),
    .A2(_0658_),
    .Y(_0693_),
    .B1(\mydesign.accum[115] ));
 sg13g2_or3_1 _3683_ (.A(_0691_),
    .B(_0692_),
    .C(_0693_),
    .X(_0694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3684_ (.B1(_0691_),
    .VDD(VPWR),
    .Y(_0695_),
    .VSS(VGND),
    .A1(_0692_),
    .A2(_0693_));
 sg13g2_and3_1 _3685_ (.X(_0696_),
    .A(_0674_),
    .B(_0694_),
    .C(_0695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3686_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0694_),
    .A2(_0695_),
    .Y(_0697_),
    .B1(_0674_));
 sg13g2_or3_1 _3687_ (.A(_0690_),
    .B(_0696_),
    .C(_0697_),
    .X(_0698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3688_ (.B1(_0690_),
    .VDD(VPWR),
    .Y(_0699_),
    .VSS(VGND),
    .A1(_0696_),
    .A2(_0697_));
 sg13g2_nand3_1 _3689_ (.B(_0698_),
    .C(_0699_),
    .A(_0678_),
    .Y(_0700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3690_ (.A2(_0699_),
    .A1(_0698_),
    .B1(_0678_),
    .X(_0701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3691_ (.X(_0702_),
    .A(_0689_),
    .B(_0700_),
    .C(_0701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3692_ (.B(_0700_),
    .C(_0701_),
    .A(_0689_),
    .Y(_0703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3693_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0700_),
    .A2(_0701_),
    .Y(_0704_),
    .B1(_0689_));
 sg13g2_nor3_1 _3694_ (.A(_0688_),
    .B(_0702_),
    .C(_0704_),
    .Y(_0705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3695_ (.B1(_0688_),
    .VDD(VPWR),
    .Y(_0706_),
    .VSS(VGND),
    .A1(_0702_),
    .A2(_0704_));
 sg13g2_nor2b_1 _3696_ (.A(_0705_),
    .B_N(_0706_),
    .Y(_0707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3697_ (.Y(_0708_),
    .A(_0687_),
    .B(_0707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3698_ (.B1(net470),
    .VDD(VPWR),
    .Y(_0709_),
    .VSS(VGND),
    .A1(net577),
    .A2(net936));
 sg13g2_a21oi_1 _3699_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net577),
    .A2(_0708_),
    .Y(_0107_),
    .B1(_0709_));
 sg13g2_nor2b_1 _3700_ (.A(_0696_),
    .B_N(_0698_),
    .Y(_0710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3701_ (.Y(_0711_),
    .A(\mydesign.pe_inputs[63] ),
    .B(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3702_ (.Y(_0712_),
    .B(_0694_),
    .A_N(_0692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3703_ (.Y(_0713_),
    .A(\mydesign.pe_inputs[62] ),
    .B(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3704_ (.A(\mydesign.pe_inputs[61] ),
    .B(_0658_),
    .X(_0714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3705_ (.Y(_0715_),
    .A(\mydesign.accum[116] ),
    .B(_0714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3706_ (.A(_0713_),
    .B(_0715_),
    .Y(_0716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3707_ (.B(_0715_),
    .A(_0713_),
    .X(_0717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3708_ (.Y(_0718_),
    .A(_0712_),
    .B(_0717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3709_ (.Y(_0719_),
    .A(_0712_),
    .B(_0717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3710_ (.B(_0719_),
    .A(_0711_),
    .X(_0720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3711_ (.Y(_0721_),
    .B(_0720_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0710_));
 sg13g2_xor2_1 _3712_ (.B(_0720_),
    .A(_0710_),
    .X(_0722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3713_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0700_),
    .A2(_0703_),
    .Y(_0723_),
    .B1(_0722_));
 sg13g2_nand3_1 _3714_ (.B(_0703_),
    .C(_0722_),
    .A(_0700_),
    .Y(_0724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3715_ (.Y(_0725_),
    .B(_0724_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0723_));
 sg13g2_a21oi_1 _3716_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0687_),
    .A2(_0706_),
    .Y(_0726_),
    .B1(_0705_));
 sg13g2_nor2_1 _3717_ (.A(_0725_),
    .B(_0726_),
    .Y(_0727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3718_ (.Y(_0728_),
    .A(_0725_),
    .B(_0726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3719_ (.B1(net470),
    .VDD(VPWR),
    .Y(_0729_),
    .VSS(VGND),
    .A1(net577),
    .A2(net972));
 sg13g2_a21oi_1 _3720_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net577),
    .A2(_0728_),
    .Y(_0108_),
    .B1(_0729_));
 sg13g2_nor2_1 _3721_ (.A(_0723_),
    .B(_0727_),
    .Y(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3722_ (.B1(_0718_),
    .VDD(VPWR),
    .Y(_0731_),
    .VSS(VGND),
    .A1(_0711_),
    .A2(_0719_));
 sg13g2_nand2_1 _3723_ (.Y(_0732_),
    .A(\mydesign.pe_inputs[63] ),
    .B(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3724_ (.B(\mydesign.pe_inputs[62] ),
    .C(_0658_),
    .A(\mydesign.accum[117] ),
    .Y(_0733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3725_ (.A2(_0658_),
    .A1(\mydesign.pe_inputs[62] ),
    .B1(\mydesign.accum[117] ),
    .X(_0734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3726_ (.Y(_0735_),
    .A(_0733_),
    .B(_0734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3727_ (.B(_0735_),
    .A(_0732_),
    .X(_0736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3728_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[116] ),
    .A2(_0714_),
    .Y(_0737_),
    .B1(_0716_));
 sg13g2_nand2b_1 _3729_ (.Y(_0738_),
    .B(_0736_),
    .A_N(_0737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3730_ (.Y(_0739_),
    .A(_0736_),
    .B(_0737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3731_ (.Y(_0740_),
    .A(_0731_),
    .B(_0739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3732_ (.Y(_0741_),
    .A(_0731_),
    .B(_0739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3733_ (.Y(_0742_),
    .A(_0721_),
    .B(_0741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3734_ (.A(_0721_),
    .B(_0741_),
    .Y(_0743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3735_ (.Y(_0744_),
    .A(_0721_),
    .B(_0741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3736_ (.Y(_0745_),
    .A(_0730_),
    .B(_0744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3737_ (.B1(net471),
    .VDD(VPWR),
    .Y(_0746_),
    .VSS(VGND),
    .A1(net580),
    .A2(net960));
 sg13g2_a21oi_1 _3738_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net577),
    .A2(_0745_),
    .Y(_0109_),
    .B1(_0746_));
 sg13g2_a21oi_1 _3739_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_inputs[63] ),
    .A2(_0658_),
    .Y(_0747_),
    .B1(\mydesign.accum[118] ));
 sg13g2_nand3_1 _3740_ (.B(\mydesign.pe_inputs[63] ),
    .C(_0658_),
    .A(\mydesign.accum[118] ),
    .Y(_0748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3741_ (.Y(_0749_),
    .B(_0748_),
    .A_N(_0747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3742_ (.B1(_0733_),
    .VDD(VPWR),
    .Y(_0750_),
    .VSS(VGND),
    .A1(_0732_),
    .A2(_0735_));
 sg13g2_inv_1 _3743_ (.VDD(VPWR),
    .Y(_0751_),
    .A(_0750_),
    .VSS(VGND));
 sg13g2_xnor2_1 _3744_ (.Y(_0752_),
    .A(_0749_),
    .B(_0750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3745_ (.Y(_0753_),
    .B(_0752_),
    .A_N(_0738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3746_ (.Y(_0754_),
    .A(_0738_),
    .B(_0752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3747_ (.Y(_0755_),
    .B(_0754_),
    .A_N(_0740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3748_ (.Y(_0756_),
    .A(_0740_),
    .B(_0754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3749_ (.A(_0723_),
    .B(_0743_),
    .Y(_0757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3750_ (.B1(_0757_),
    .VDD(VPWR),
    .Y(_0758_),
    .VSS(VGND),
    .A1(_0725_),
    .A2(_0726_));
 sg13g2_a21o_1 _3751_ (.A2(_0758_),
    .A1(_0742_),
    .B1(_0756_),
    .X(_0759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3752_ (.B(_0756_),
    .C(_0758_),
    .A(_0742_),
    .Y(_0760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3753_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0759_),
    .A2(_0760_),
    .Y(_0761_),
    .B1(net502));
 sg13g2_o21ai_1 _3754_ (.B1(net471),
    .VDD(VPWR),
    .Y(_0762_),
    .VSS(VGND),
    .A1(net570),
    .A2(net898));
 sg13g2_nor2_1 _3755_ (.A(_0761_),
    .B(_0762_),
    .Y(_0110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3756_ (.Y(_0763_),
    .A(_0755_),
    .B(_0760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3757_ (.B1(_0748_),
    .VDD(VPWR),
    .Y(_0764_),
    .VSS(VGND),
    .A1(_0747_),
    .A2(_0751_));
 sg13g2_xor2_1 _3758_ (.B(_0764_),
    .A(net973),
    .X(_0765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3759_ (.Y(_0766_),
    .A(_0753_),
    .B(_0765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3760_ (.Y(_0767_),
    .A(_0763_),
    .B(_0766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3761_ (.B1(net471),
    .VDD(VPWR),
    .Y(_0768_),
    .VSS(VGND),
    .A1(net571),
    .A2(net973));
 sg13g2_a21oi_1 _3762_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net570),
    .A2(_0767_),
    .Y(_0111_),
    .B1(_0768_));
 sg13g2_nand3_1 _3763_ (.B(_2638_),
    .C(_2647_),
    .A(net610),
    .Y(_0769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3764_ (.A(net612),
    .B(_0769_),
    .X(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3765_ (.Y(_0771_),
    .A(net411),
    .B(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3766_ (.B1(_0771_),
    .VDD(VPWR),
    .Y(_0112_),
    .VSS(VGND),
    .A1(net603),
    .A2(_0769_));
 sg13g2_nand2_1 _3767_ (.Y(_0772_),
    .A(net672),
    .B(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3768_ (.B1(_0772_),
    .VDD(VPWR),
    .Y(_0113_),
    .VSS(VGND),
    .A1(net601),
    .A2(_0769_));
 sg13g2_nand2_1 _3769_ (.Y(_0773_),
    .A(net701),
    .B(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3770_ (.B1(_0773_),
    .VDD(VPWR),
    .Y(_0114_),
    .VSS(VGND),
    .A1(net599),
    .A2(_0769_));
 sg13g2_nand2_1 _3771_ (.Y(_0774_),
    .A(net707),
    .B(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3772_ (.B1(_0774_),
    .VDD(VPWR),
    .Y(_0115_),
    .VSS(VGND),
    .A1(net597),
    .A2(_0769_));
 sg13g2_o21ai_1 _3773_ (.B1(net622),
    .VDD(VPWR),
    .Y(_0775_),
    .VSS(VGND),
    .A1(net1076),
    .A2(net433));
 sg13g2_a21oi_1 _3774_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2583_),
    .A2(net433),
    .Y(_0116_),
    .B1(_0775_));
 sg13g2_o21ai_1 _3775_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0776_),
    .VSS(VGND),
    .A1(net1024),
    .A2(net433));
 sg13g2_a21oi_1 _3776_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2582_),
    .A2(net433),
    .Y(_0117_),
    .B1(_0776_));
 sg13g2_o21ai_1 _3777_ (.B1(net627),
    .VDD(VPWR),
    .Y(_0777_),
    .VSS(VGND),
    .A1(net1036),
    .A2(net433));
 sg13g2_a21oi_1 _3778_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2581_),
    .A2(net435),
    .Y(_0118_),
    .B1(_0777_));
 sg13g2_o21ai_1 _3779_ (.B1(net622),
    .VDD(VPWR),
    .Y(_0778_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[55] ),
    .A2(net435));
 sg13g2_a21oi_1 _3780_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2580_),
    .A2(net435),
    .Y(_0119_),
    .B1(_0778_));
 sg13g2_a21oi_1 _3781_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net497),
    .A2(_2589_),
    .Y(_0779_),
    .B1(_0393_));
 sg13g2_o21ai_1 _3782_ (.B1(_0779_),
    .VDD(VPWR),
    .Y(_0780_),
    .VSS(VGND),
    .A1(net497),
    .A2(\mydesign.weights[2][12] ));
 sg13g2_nor2_1 _3783_ (.A(net497),
    .B(\mydesign.weights[2][4] ),
    .Y(_0781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3784_ (.B1(net459),
    .VDD(VPWR),
    .Y(_0782_),
    .VSS(VGND),
    .A1(net552),
    .A2(\mydesign.weights[2][8] ));
 sg13g2_o21ai_1 _3785_ (.B1(_0780_),
    .VDD(VPWR),
    .Y(_0783_),
    .VSS(VGND),
    .A1(_0781_),
    .A2(_0782_));
 sg13g2_o21ai_1 _3786_ (.B1(net629),
    .VDD(VPWR),
    .Y(_0784_),
    .VSS(VGND),
    .A1(net491),
    .A2(_0783_));
 sg13g2_a21oi_1 _3787_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2559_),
    .A2(net491),
    .Y(_0120_),
    .B1(_0784_));
 sg13g2_nor2_1 _3788_ (.A(net497),
    .B(\mydesign.weights[2][5] ),
    .Y(_0785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3789_ (.B1(net459),
    .VDD(VPWR),
    .Y(_0786_),
    .VSS(VGND),
    .A1(net550),
    .A2(\mydesign.weights[2][9] ));
 sg13g2_mux2_1 _3790_ (.A0(\mydesign.weights[2][17] ),
    .A1(\mydesign.weights[2][13] ),
    .S(net551),
    .X(_0787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3791_ (.Y(_0788_),
    .A(_0392_),
    .B(_0787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3792_ (.B1(_0788_),
    .VDD(VPWR),
    .Y(_0789_),
    .VSS(VGND),
    .A1(_0785_),
    .A2(_0786_));
 sg13g2_o21ai_1 _3793_ (.B1(net629),
    .VDD(VPWR),
    .Y(_0790_),
    .VSS(VGND),
    .A1(net491),
    .A2(_0789_));
 sg13g2_a21oi_1 _3794_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2558_),
    .A2(net491),
    .Y(_0121_),
    .B1(_0790_));
 sg13g2_nand2b_1 _3795_ (.Y(_0791_),
    .B(net551),
    .A_N(\mydesign.weights[2][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3796_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0792_),
    .B(\mydesign.weights[2][10] ),
    .A(net549));
 sg13g2_nand3_1 _3797_ (.B(_0791_),
    .C(_0792_),
    .A(net459),
    .Y(_0793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3798_ (.A0(\mydesign.weights[2][18] ),
    .A1(\mydesign.weights[2][14] ),
    .S(net551),
    .X(_0794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3799_ (.Y(_0795_),
    .A(_0392_),
    .B(_0794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3800_ (.Y(_0796_),
    .A(_0793_),
    .B(_0795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3801_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0797_),
    .VSS(VGND),
    .A1(net491),
    .A2(_0796_));
 sg13g2_a21oi_1 _3802_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2557_),
    .A2(net491),
    .Y(_0122_),
    .B1(_0797_));
 sg13g2_nor2b_1 _3803_ (.A(\mydesign.weights[2][7] ),
    .B_N(net551),
    .Y(_0798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3804_ (.A(net550),
    .B(\mydesign.weights[2][11] ),
    .Y(_0799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3805_ (.A(_0397_),
    .B(_0798_),
    .C(_0799_),
    .Y(_0800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3806_ (.A(net550),
    .B(\mydesign.weights[2][19] ),
    .Y(_0801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3807_ (.A(\mydesign.weights[2][15] ),
    .B_N(net550),
    .Y(_0802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3808_ (.A(_0393_),
    .B(_0801_),
    .C(_0802_),
    .Y(_0803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3809_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0804_),
    .B(_0803_),
    .A(_0800_));
 sg13g2_o21ai_1 _3810_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0805_),
    .VSS(VGND),
    .A1(net491),
    .A2(_0804_));
 sg13g2_a21oi_1 _3811_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2556_),
    .A2(net492),
    .Y(_0123_),
    .B1(_0805_));
 sg13g2_and3_1 _3812_ (.X(_0806_),
    .A(net572),
    .B(\mydesign.pe_inputs[56] ),
    .C(_0783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3813_ (.B1(net474),
    .VDD(VPWR),
    .Y(_0807_),
    .VSS(VGND),
    .A1(net688),
    .A2(_0806_));
 sg13g2_a21oi_1 _3814_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net688),
    .A2(_0806_),
    .Y(_0124_),
    .B1(_0807_));
 sg13g2_nand3_1 _3815_ (.B(\mydesign.pe_inputs[56] ),
    .C(_0789_),
    .A(\mydesign.accum[105] ),
    .Y(_0808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3816_ (.A2(_0789_),
    .A1(\mydesign.pe_inputs[56] ),
    .B1(\mydesign.accum[105] ),
    .X(_0809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3817_ (.Y(_0810_),
    .A(_0808_),
    .B(_0809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3818_ (.Y(_0811_),
    .A(\mydesign.pe_inputs[57] ),
    .B(_0783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3819_ (.A(_0810_),
    .B(_0811_),
    .Y(_0812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3820_ (.B(_0811_),
    .A(_0810_),
    .X(_0813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3821_ (.B(\mydesign.pe_inputs[56] ),
    .C(_0783_),
    .A(net688),
    .Y(_0814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3822_ (.B(\mydesign.pe_inputs[56] ),
    .C(_0783_),
    .A(net688),
    .Y(_0815_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0813_));
 sg13g2_xor2_1 _3823_ (.B(_0814_),
    .A(_0813_),
    .X(_0816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3824_ (.B1(net465),
    .VDD(VPWR),
    .Y(_0817_),
    .VSS(VGND),
    .A1(net572),
    .A2(net916));
 sg13g2_a21oi_1 _3825_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net572),
    .A2(_0816_),
    .Y(_0125_),
    .B1(_0817_));
 sg13g2_nand2_1 _3826_ (.Y(_0818_),
    .A(\mydesign.pe_inputs[58] ),
    .B(_0783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3827_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0793_),
    .A2(_0795_),
    .Y(_0819_),
    .B1(_2583_));
 sg13g2_nand2_1 _3828_ (.Y(_0820_),
    .A(\mydesign.accum[106] ),
    .B(_0819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3829_ (.B(_0819_),
    .A(\mydesign.accum[106] ),
    .X(_0821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3830_ (.Y(_0822_),
    .A(\mydesign.pe_inputs[57] ),
    .B(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3831_ (.X(_0823_),
    .A(\mydesign.pe_inputs[57] ),
    .B(_0789_),
    .C(_0821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3832_ (.Y(_0824_),
    .A(_0821_),
    .B(_0822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3833_ (.VDD(VPWR),
    .Y(_0825_),
    .A(_0824_),
    .VSS(VGND));
 sg13g2_xnor2_1 _3834_ (.Y(_0826_),
    .A(_0808_),
    .B(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3835_ (.Y(_0827_),
    .B(_0826_),
    .A_N(_0818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3836_ (.Y(_0828_),
    .A(_0818_),
    .B(_0826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3837_ (.Y(_0829_),
    .A(_0812_),
    .B(_0828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3838_ (.Y(_0830_),
    .A(_0812_),
    .B(_0828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3839_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0831_),
    .B(_0830_),
    .A(_0815_));
 sg13g2_xnor2_1 _3840_ (.Y(_0832_),
    .A(_0815_),
    .B(_0830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3841_ (.B1(net465),
    .VDD(VPWR),
    .Y(_0833_),
    .VSS(VGND),
    .A1(net572),
    .A2(net1010));
 sg13g2_a21oi_1 _3842_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net572),
    .A2(_0832_),
    .Y(_0126_),
    .B1(_0833_));
 sg13g2_and2_1 _3843_ (.A(_0829_),
    .B(_0831_),
    .X(_0834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3844_ (.B1(_0827_),
    .VDD(VPWR),
    .Y(_0835_),
    .VSS(VGND),
    .A1(_0808_),
    .A2(_0825_));
 sg13g2_nand2_1 _3845_ (.Y(_0836_),
    .A(\mydesign.pe_inputs[59] ),
    .B(_0783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3846_ (.Y(_0837_),
    .A(\mydesign.pe_inputs[58] ),
    .B(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3847_ (.Y(_0838_),
    .A(\mydesign.pe_inputs[57] ),
    .B(_0796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3848_ (.B1(\mydesign.pe_inputs[56] ),
    .VDD(VPWR),
    .Y(_0839_),
    .VSS(VGND),
    .A1(_0800_),
    .A2(_0803_));
 sg13g2_nand3_1 _3849_ (.B(\mydesign.pe_inputs[56] ),
    .C(_0804_),
    .A(\mydesign.accum[107] ),
    .Y(_0840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3850_ (.B(_0839_),
    .A(\mydesign.accum[107] ),
    .X(_0841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3851_ (.B(_0841_),
    .A(_0838_),
    .X(_0842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3852_ (.VDD(VPWR),
    .Y(_0843_),
    .A(_0842_),
    .VSS(VGND));
 sg13g2_xnor2_1 _3853_ (.Y(_0844_),
    .A(_0820_),
    .B(_0842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3854_ (.Y(_0845_),
    .B(_0844_),
    .A_N(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3855_ (.Y(_0846_),
    .A(_0837_),
    .B(_0844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3856_ (.Y(_0847_),
    .A(_0823_),
    .B(_0846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3857_ (.A(_0823_),
    .B(_0846_),
    .Y(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3858_ (.B(_0846_),
    .A(_0823_),
    .X(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3859_ (.Y(_0850_),
    .A(_0836_),
    .B(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3860_ (.Y(_0851_),
    .A(_0835_),
    .B(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3861_ (.Y(_0852_),
    .A(_0835_),
    .B(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3862_ (.Y(_0853_),
    .A(_0834_),
    .B(_0852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3863_ (.B1(net465),
    .VDD(VPWR),
    .Y(_0854_),
    .VSS(VGND),
    .A1(net572),
    .A2(net1009));
 sg13g2_a21oi_1 _3864_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net572),
    .A2(_0853_),
    .Y(_0127_),
    .B1(_0854_));
 sg13g2_o21ai_1 _3865_ (.B1(_0851_),
    .VDD(VPWR),
    .Y(_0855_),
    .VSS(VGND),
    .A1(_0834_),
    .A2(_0852_));
 sg13g2_o21ai_1 _3866_ (.B1(_0845_),
    .VDD(VPWR),
    .Y(_0856_),
    .VSS(VGND),
    .A1(_0820_),
    .A2(_0843_));
 sg13g2_nand2_1 _3867_ (.Y(_0857_),
    .A(\mydesign.pe_inputs[59] ),
    .B(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3868_ (.B1(_0840_),
    .VDD(VPWR),
    .Y(_0858_),
    .VSS(VGND),
    .A1(_0838_),
    .A2(_0841_));
 sg13g2_nand2_1 _3869_ (.Y(_0859_),
    .A(\mydesign.pe_inputs[58] ),
    .B(_0796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3870_ (.B(\mydesign.pe_inputs[57] ),
    .C(_0804_),
    .A(\mydesign.accum[108] ),
    .Y(_0860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3871_ (.A2(_0804_),
    .A1(\mydesign.pe_inputs[57] ),
    .B1(\mydesign.accum[108] ),
    .X(_0861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3872_ (.Y(_0862_),
    .A(_0860_),
    .B(_0861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3873_ (.B(_0862_),
    .A(_0859_),
    .X(_0863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3874_ (.A(_0858_),
    .B(_0863_),
    .X(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3875_ (.Y(_0865_),
    .A(_0858_),
    .B(_0863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3876_ (.A(_0857_),
    .B(_0865_),
    .Y(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3877_ (.B(_0865_),
    .A(_0857_),
    .X(_0867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3878_ (.Y(_0868_),
    .A(_0856_),
    .B(_0867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3879_ (.Y(_0869_),
    .A(_0856_),
    .B(_0867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3880_ (.B1(_0847_),
    .VDD(VPWR),
    .Y(_0870_),
    .VSS(VGND),
    .A1(_0836_),
    .A2(_0848_));
 sg13g2_nor2b_1 _3881_ (.A(_0869_),
    .B_N(_0870_),
    .Y(_0871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3882_ (.Y(_0872_),
    .B(_0869_),
    .A_N(_0870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3883_ (.Y(_0873_),
    .B(_0872_),
    .A_N(_0871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3884_ (.Y(_0874_),
    .A(_0855_),
    .B(_0873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3885_ (.B1(net465),
    .VDD(VPWR),
    .Y(_0875_),
    .VSS(VGND),
    .A1(net501),
    .A2(_0874_));
 sg13g2_a21oi_1 _3886_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net501),
    .A2(_2579_),
    .Y(_0128_),
    .B1(_0875_));
 sg13g2_a21oi_1 _3887_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0855_),
    .A2(_0872_),
    .Y(_0876_),
    .B1(_0871_));
 sg13g2_nand2_1 _3888_ (.Y(_0877_),
    .A(\mydesign.pe_inputs[59] ),
    .B(_0796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3889_ (.A(\mydesign.pe_inputs[58] ),
    .B(_0804_),
    .X(_0878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3890_ (.Y(_0879_),
    .A(\mydesign.accum[109] ),
    .B(_0878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3891_ (.A(_0877_),
    .B(_0879_),
    .Y(_0880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3892_ (.B(_0879_),
    .A(_0877_),
    .X(_0881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3893_ (.B1(_0860_),
    .VDD(VPWR),
    .Y(_0882_),
    .VSS(VGND),
    .A1(_0859_),
    .A2(_0862_));
 sg13g2_nand2_1 _3894_ (.Y(_0883_),
    .A(_0881_),
    .B(_0882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3895_ (.B(_0882_),
    .A(_0881_),
    .X(_0884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3896_ (.B1(_0884_),
    .VDD(VPWR),
    .Y(_0885_),
    .VSS(VGND),
    .A1(_0864_),
    .A2(_0866_));
 sg13g2_or3_1 _3897_ (.A(_0864_),
    .B(_0866_),
    .C(_0884_),
    .X(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3898_ (.Y(_0887_),
    .A(_0885_),
    .B(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3899_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0888_),
    .B(_0887_),
    .A(_0868_));
 sg13g2_xnor2_1 _3900_ (.Y(_0889_),
    .A(_0868_),
    .B(_0887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3901_ (.Y(_0890_),
    .A(_0876_),
    .B(_0889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3902_ (.B1(net465),
    .VDD(VPWR),
    .Y(_0891_),
    .VSS(VGND),
    .A1(net573),
    .A2(net942));
 sg13g2_a21oi_1 _3903_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net572),
    .A2(_0890_),
    .Y(_0129_),
    .B1(_0891_));
 sg13g2_o21ai_1 _3904_ (.B1(_0888_),
    .VDD(VPWR),
    .Y(_0892_),
    .VSS(VGND),
    .A1(_0876_),
    .A2(_0889_));
 sg13g2_a21oi_1 _3905_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_inputs[59] ),
    .A2(_0804_),
    .Y(_0893_),
    .B1(\mydesign.accum[110] ));
 sg13g2_nand3_1 _3906_ (.B(\mydesign.pe_inputs[59] ),
    .C(_0804_),
    .A(\mydesign.accum[110] ),
    .Y(_0894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3907_ (.Y(_0895_),
    .B(_0894_),
    .A_N(_0893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3908_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[109] ),
    .A2(_0878_),
    .Y(_0896_),
    .B1(_0880_));
 sg13g2_xnor2_1 _3909_ (.Y(_0897_),
    .A(_0895_),
    .B(_0896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3910_ (.A(_0883_),
    .B(_0897_),
    .Y(_0898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3911_ (.B(_0897_),
    .A(_0883_),
    .X(_0899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3912_ (.A(_0885_),
    .B_N(_0899_),
    .Y(_0900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3913_ (.Y(_0901_),
    .A(_0885_),
    .B(_0899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3914_ (.Y(_0902_),
    .A(_0892_),
    .B(_0901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3915_ (.B1(net470),
    .VDD(VPWR),
    .Y(_0903_),
    .VSS(VGND),
    .A1(net570),
    .A2(net998));
 sg13g2_a21oi_1 _3916_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net570),
    .A2(_0902_),
    .Y(_0130_),
    .B1(_0903_));
 sg13g2_a21oi_1 _3917_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0892_),
    .A2(_0901_),
    .Y(_0904_),
    .B1(_0900_));
 sg13g2_o21ai_1 _3918_ (.B1(_0894_),
    .VDD(VPWR),
    .Y(_0905_),
    .VSS(VGND),
    .A1(_0893_),
    .A2(_0896_));
 sg13g2_xnor2_1 _3919_ (.Y(_0906_),
    .A(net835),
    .B(_0905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3920_ (.B(_0906_),
    .A(_0898_),
    .X(_0907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3921_ (.Y(_0908_),
    .A(_0904_),
    .B(_0907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3922_ (.B1(net472),
    .VDD(VPWR),
    .Y(_0909_),
    .VSS(VGND),
    .A1(net578),
    .A2(net835));
 sg13g2_a21oi_1 _3923_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net578),
    .A2(_0908_),
    .Y(_0131_),
    .B1(_0909_));
 sg13g2_o21ai_1 _3924_ (.B1(net615),
    .VDD(VPWR),
    .Y(_0910_),
    .VSS(VGND),
    .A1(_2622_),
    .A2(_2683_));
 sg13g2_nand2_2 _3925_ (.Y(_0911_),
    .A(_2655_),
    .B(_0910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3926_ (.A0(_2667_),
    .A1(net783),
    .S(_0911_),
    .X(_0132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3927_ (.A0(_2668_),
    .A1(net768),
    .S(_0911_),
    .X(_0133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3928_ (.A0(_2669_),
    .A1(net785),
    .S(_0911_),
    .X(_0134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3929_ (.A0(_2670_),
    .A1(net792),
    .S(_0911_),
    .X(_0135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3930_ (.B1(net459),
    .VDD(VPWR),
    .Y(_0912_),
    .VSS(VGND),
    .A1(\mydesign.weights[3][8] ),
    .A2(net547));
 sg13g2_a21oi_1 _3931_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net547),
    .A2(_2593_),
    .Y(_0913_),
    .B1(_0912_));
 sg13g2_a221oi_1 _3932_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net985),
    .C1(_0913_),
    .B1(_0395_),
    .A1(net725),
    .Y(_0914_),
    .A2(net454));
 sg13g2_o21ai_1 _3933_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0915_),
    .VSS(VGND),
    .A1(net1091),
    .A2(net433));
 sg13g2_a21oi_1 _3934_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net433),
    .A2(_0914_),
    .Y(_0136_),
    .B1(_0915_));
 sg13g2_nor2_1 _3935_ (.A(net497),
    .B(\mydesign.weights[3][5] ),
    .Y(_0916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3936_ (.B1(net459),
    .VDD(VPWR),
    .Y(_0917_),
    .VSS(VGND),
    .A1(\mydesign.weights[3][9] ),
    .A2(net547));
 sg13g2_a22oi_1 _3937_ (.Y(_0918_),
    .B1(_0395_),
    .B2(\mydesign.weights[3][13] ),
    .A2(net454),
    .A1(\mydesign.weights[3][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3938_ (.B1(_0918_),
    .VDD(VPWR),
    .Y(_0919_),
    .VSS(VGND),
    .A1(_0916_),
    .A2(_0917_));
 sg13g2_o21ai_1 _3939_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0920_),
    .VSS(VGND),
    .A1(net486),
    .A2(_0919_));
 sg13g2_a21oi_1 _3940_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2555_),
    .A2(net486),
    .Y(_0137_),
    .B1(_0920_));
 sg13g2_nand2b_1 _3941_ (.Y(_0921_),
    .B(\mydesign.weights[3][10] ),
    .A_N(net547),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3942_ (.Y(_0922_),
    .A(net547),
    .B(\mydesign.weights[3][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3943_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0921_),
    .A2(_0922_),
    .Y(_0923_),
    .B1(_0397_));
 sg13g2_and3_1 _3944_ (.X(_0924_),
    .A(net541),
    .B(\mydesign.weights[3][2] ),
    .C(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3945_ (.X(_0925_),
    .A(\mydesign.weights[3][14] ),
    .B(net547),
    .C(_0392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3946_ (.A(_0923_),
    .B(_0924_),
    .C(_0925_),
    .X(_0926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3947_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0927_),
    .VSS(VGND),
    .A1(net486),
    .A2(_0926_));
 sg13g2_a21oi_1 _3948_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2554_),
    .A2(net486),
    .Y(_0138_),
    .B1(_0927_));
 sg13g2_nand2b_1 _3949_ (.Y(_0928_),
    .B(\mydesign.weights[3][11] ),
    .A_N(net548),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3950_ (.Y(_0929_),
    .A(net547),
    .B(\mydesign.weights[3][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3951_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0928_),
    .A2(_0929_),
    .Y(_0930_),
    .B1(_0397_));
 sg13g2_and3_1 _3952_ (.X(_0931_),
    .A(\mydesign.weights[3][15] ),
    .B(_2586_),
    .C(_0394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3953_ (.X(_0932_),
    .A(net541),
    .B(\mydesign.weights[3][3] ),
    .C(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3954_ (.A(_0930_),
    .B(_0931_),
    .C(_0932_),
    .X(_0933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3955_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0934_),
    .VSS(VGND),
    .A1(net486),
    .A2(net428));
 sg13g2_a21oi_1 _3956_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2553_),
    .A2(net486),
    .Y(_0139_),
    .B1(_0934_));
 sg13g2_nor2b_1 _3957_ (.A(_0914_),
    .B_N(\mydesign.pe_inputs[52] ),
    .Y(_0935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3958_ (.Y(_0936_),
    .A(net564),
    .B(_0935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3959_ (.B(_0936_),
    .A(net1053),
    .X(_0937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3960_ (.A(net462),
    .B(net1054),
    .Y(_0140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3961_ (.B(\mydesign.pe_inputs[52] ),
    .C(_0919_),
    .A(\mydesign.accum[97] ),
    .Y(_0938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3962_ (.VDD(VPWR),
    .Y(_0939_),
    .A(_0938_),
    .VSS(VGND));
 sg13g2_a21oi_1 _3963_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_inputs[52] ),
    .A2(_0919_),
    .Y(_0940_),
    .B1(\mydesign.accum[97] ));
 sg13g2_or2_1 _3964_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0941_),
    .B(_0940_),
    .A(_0939_));
 sg13g2_nor2b_1 _3965_ (.A(_0914_),
    .B_N(\mydesign.pe_inputs[53] ),
    .Y(_0942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3966_ (.A(_0941_),
    .B_N(_0942_),
    .Y(_0943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3967_ (.Y(_0944_),
    .A(_0941_),
    .B(_0942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3968_ (.B(_0935_),
    .C(_0944_),
    .A(\mydesign.accum[96] ),
    .Y(_0945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3969_ (.A2(_0935_),
    .A1(\mydesign.accum[96] ),
    .B1(_0944_),
    .X(_0946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3970_ (.Y(_0947_),
    .A(_0945_),
    .B(_0946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3971_ (.B1(net464),
    .VDD(VPWR),
    .Y(_0948_),
    .VSS(VGND),
    .A1(net564),
    .A2(net1007));
 sg13g2_a21oi_1 _3972_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net564),
    .A2(_0947_),
    .Y(_0141_),
    .B1(_0948_));
 sg13g2_nand2b_1 _3973_ (.Y(_0949_),
    .B(\mydesign.pe_inputs[54] ),
    .A_N(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3974_ (.B(\mydesign.pe_inputs[52] ),
    .C(_0926_),
    .A(\mydesign.accum[98] ),
    .Y(_0950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3975_ (.VDD(VPWR),
    .Y(_0951_),
    .A(_0950_),
    .VSS(VGND));
 sg13g2_a21o_1 _3976_ (.A2(_0926_),
    .A1(\mydesign.pe_inputs[52] ),
    .B1(\mydesign.accum[98] ),
    .X(_0952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3977_ (.A(\mydesign.pe_inputs[53] ),
    .B(_0919_),
    .C(_0950_),
    .D(_0952_),
    .X(_0953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3978_ (.Y(_0954_),
    .B1(_0950_),
    .B2(_0952_),
    .A2(_0919_),
    .A1(\mydesign.pe_inputs[53] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3979_ (.A(_0953_),
    .B(_0954_),
    .Y(_0955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3980_ (.Y(_0956_),
    .A(_0938_),
    .B(_0955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3981_ (.A(_0949_),
    .B_N(_0956_),
    .Y(_0957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3982_ (.Y(_0958_),
    .A(_0949_),
    .B(_0956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3983_ (.Y(_0959_),
    .A(_0943_),
    .B(_0958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3984_ (.Y(_0960_),
    .A(_0943_),
    .B(_0958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3985_ (.Y(_0961_),
    .A(_0945_),
    .B(_0960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3986_ (.B1(net464),
    .VDD(VPWR),
    .Y(_0962_),
    .VSS(VGND),
    .A1(net565),
    .A2(net847));
 sg13g2_a21oi_1 _3987_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net564),
    .A2(_0961_),
    .Y(_0142_),
    .B1(_0962_));
 sg13g2_o21ai_1 _3988_ (.B1(_0959_),
    .VDD(VPWR),
    .Y(_0963_),
    .VSS(VGND),
    .A1(_0945_),
    .A2(_0960_));
 sg13g2_a21oi_1 _3989_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0939_),
    .A2(_0955_),
    .Y(_0964_),
    .B1(_0957_));
 sg13g2_nand2b_1 _3990_ (.Y(_0965_),
    .B(\mydesign.pe_inputs[55] ),
    .A_N(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3991_ (.VDD(VPWR),
    .Y(_0966_),
    .A(_0965_),
    .VSS(VGND));
 sg13g2_nand2_1 _3992_ (.Y(_0967_),
    .A(\mydesign.pe_inputs[54] ),
    .B(_0919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3993_ (.Y(_0968_),
    .A(\mydesign.pe_inputs[53] ),
    .B(_0926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3994_ (.X(_0969_),
    .A(\mydesign.accum[99] ),
    .B(\mydesign.pe_inputs[52] ),
    .C(net428),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3995_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_inputs[52] ),
    .A2(net428),
    .Y(_0970_),
    .B1(\mydesign.accum[99] ));
 sg13g2_or3_1 _3996_ (.A(_0968_),
    .B(_0969_),
    .C(_0970_),
    .X(_0971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3997_ (.B1(_0968_),
    .VDD(VPWR),
    .Y(_0972_),
    .VSS(VGND),
    .A1(_0969_),
    .A2(_0970_));
 sg13g2_and3_1 _3998_ (.X(_0973_),
    .A(_0951_),
    .B(_0971_),
    .C(_0972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3999_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0971_),
    .A2(_0972_),
    .Y(_0974_),
    .B1(_0951_));
 sg13g2_or3_1 _4000_ (.A(_0967_),
    .B(_0973_),
    .C(_0974_),
    .X(_0975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4001_ (.B1(_0967_),
    .VDD(VPWR),
    .Y(_0976_),
    .VSS(VGND),
    .A1(_0973_),
    .A2(_0974_));
 sg13g2_and2_1 _4002_ (.A(_0975_),
    .B(_0976_),
    .X(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4003_ (.B(_0975_),
    .C(_0976_),
    .A(_0953_),
    .Y(_0978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4004_ (.A2(_0976_),
    .A1(_0975_),
    .B1(_0953_),
    .X(_0979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4005_ (.X(_0980_),
    .A(_0966_),
    .B(_0978_),
    .C(_0979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4006_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0978_),
    .A2(_0979_),
    .Y(_0981_),
    .B1(_0966_));
 sg13g2_nor3_1 _4007_ (.A(_0964_),
    .B(_0980_),
    .C(_0981_),
    .Y(_0982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4008_ (.B1(_0964_),
    .VDD(VPWR),
    .Y(_0983_),
    .VSS(VGND),
    .A1(_0980_),
    .A2(_0981_));
 sg13g2_nor2b_1 _4009_ (.A(_0982_),
    .B_N(_0983_),
    .Y(_0984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4010_ (.Y(_0985_),
    .A(_0963_),
    .B(_0984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4011_ (.B1(net466),
    .VDD(VPWR),
    .Y(_0986_),
    .VSS(VGND),
    .A1(net564),
    .A2(net967));
 sg13g2_a21oi_1 _4012_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net564),
    .A2(_0985_),
    .Y(_0143_),
    .B1(_0986_));
 sg13g2_nor2b_1 _4013_ (.A(_0973_),
    .B_N(_0975_),
    .Y(_0987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4014_ (.Y(_0988_),
    .A(\mydesign.pe_inputs[55] ),
    .B(_0919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4015_ (.Y(_0989_),
    .B(_0971_),
    .A_N(_0969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4016_ (.Y(_0990_),
    .A(\mydesign.pe_inputs[54] ),
    .B(_0926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4017_ (.B(\mydesign.pe_inputs[53] ),
    .C(net428),
    .A(\mydesign.accum[100] ),
    .Y(_0991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4018_ (.A2(_0933_),
    .A1(\mydesign.pe_inputs[53] ),
    .B1(\mydesign.accum[100] ),
    .X(_0992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4019_ (.Y(_0993_),
    .A(_0991_),
    .B(_0992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4020_ (.B(_0993_),
    .A(_0990_),
    .X(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4021_ (.Y(_0995_),
    .A(_0989_),
    .B(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4022_ (.Y(_0996_),
    .A(_0989_),
    .B(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4023_ (.B(_0996_),
    .A(_0988_),
    .X(_0997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4024_ (.Y(_0998_),
    .B(_0997_),
    .A_N(_0987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4025_ (.Y(_0999_),
    .A(_0987_),
    .B(_0997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4026_ (.A2(_0977_),
    .A1(_0953_),
    .B1(_0980_),
    .X(_1000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4027_ (.Y(_1001_),
    .A(_0999_),
    .B(_1000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4028_ (.B(_1000_),
    .A(_0999_),
    .X(_1002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4029_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0963_),
    .A2(_0983_),
    .Y(_1003_),
    .B1(_0982_));
 sg13g2_nand2b_1 _4030_ (.Y(_1004_),
    .B(_1002_),
    .A_N(_1003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4031_ (.B(_1003_),
    .A(_1002_),
    .X(_1005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4032_ (.B1(net466),
    .VDD(VPWR),
    .Y(_1006_),
    .VSS(VGND),
    .A1(net564),
    .A2(net1006));
 sg13g2_a21oi_1 _4033_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net564),
    .A2(_1005_),
    .Y(_0144_),
    .B1(_1006_));
 sg13g2_nand2_1 _4034_ (.Y(_1007_),
    .A(_1001_),
    .B(_1004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4035_ (.B1(_0995_),
    .VDD(VPWR),
    .Y(_1008_),
    .VSS(VGND),
    .A1(_0988_),
    .A2(_0996_));
 sg13g2_nand2_1 _4036_ (.Y(_1009_),
    .A(\mydesign.pe_inputs[55] ),
    .B(_0926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4037_ (.B(\mydesign.pe_inputs[54] ),
    .C(net428),
    .A(\mydesign.accum[101] ),
    .Y(_1010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4038_ (.A2(net428),
    .A1(\mydesign.pe_inputs[54] ),
    .B1(\mydesign.accum[101] ),
    .X(_1011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4039_ (.Y(_1012_),
    .A(_1010_),
    .B(_1011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4040_ (.B(_1012_),
    .A(_1009_),
    .X(_1013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4041_ (.B1(_0991_),
    .VDD(VPWR),
    .Y(_1014_),
    .VSS(VGND),
    .A1(_0990_),
    .A2(_0993_));
 sg13g2_nand2_1 _4042_ (.Y(_1015_),
    .A(_1013_),
    .B(_1014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4043_ (.B(_1014_),
    .A(_1013_),
    .X(_1016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4044_ (.Y(_1017_),
    .A(_1008_),
    .B(_1016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4045_ (.Y(_1018_),
    .A(_1008_),
    .B(_1016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4046_ (.Y(_1019_),
    .A(_0998_),
    .B(_1018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4047_ (.B(_1019_),
    .A(_1007_),
    .X(_1020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4048_ (.B1(net464),
    .VDD(VPWR),
    .Y(_1021_),
    .VSS(VGND),
    .A1(net565),
    .A2(net968));
 sg13g2_a21oi_1 _4049_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net565),
    .A2(_1020_),
    .Y(_0145_),
    .B1(_1021_));
 sg13g2_a21o_1 _4050_ (.A2(_1001_),
    .A1(_0998_),
    .B1(_1018_),
    .X(_1022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4051_ (.B1(_1022_),
    .VDD(VPWR),
    .Y(_1023_),
    .VSS(VGND),
    .A1(_1004_),
    .A2(_1019_));
 sg13g2_a21oi_1 _4052_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_inputs[55] ),
    .A2(net428),
    .Y(_1024_),
    .B1(\mydesign.accum[102] ));
 sg13g2_nand3_1 _4053_ (.B(\mydesign.pe_inputs[55] ),
    .C(net428),
    .A(\mydesign.accum[102] ),
    .Y(_1025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4054_ (.Y(_1026_),
    .B(_1025_),
    .A_N(_1024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4055_ (.B1(_1010_),
    .VDD(VPWR),
    .Y(_1027_),
    .VSS(VGND),
    .A1(_1009_),
    .A2(_1012_));
 sg13g2_inv_1 _4056_ (.VDD(VPWR),
    .Y(_1028_),
    .A(_1027_),
    .VSS(VGND));
 sg13g2_xnor2_1 _4057_ (.Y(_1029_),
    .A(_1026_),
    .B(_1027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4058_ (.Y(_1030_),
    .B(_1029_),
    .A_N(_1015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4059_ (.Y(_1031_),
    .A(_1015_),
    .B(_1029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4060_ (.B(_1016_),
    .C(_1031_),
    .A(_1008_),
    .Y(_1032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4061_ (.VDD(VPWR),
    .Y(_1033_),
    .A(_1032_),
    .VSS(VGND));
 sg13g2_xnor2_1 _4062_ (.Y(_1034_),
    .A(_1017_),
    .B(_1031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4063_ (.Y(_1035_),
    .A(_1023_),
    .B(_1034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4064_ (.B1(net464),
    .VDD(VPWR),
    .Y(_1036_),
    .VSS(VGND),
    .A1(net566),
    .A2(net944));
 sg13g2_a21oi_1 _4065_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net566),
    .A2(_1035_),
    .Y(_0146_),
    .B1(_1036_));
 sg13g2_a21oi_1 _4066_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1023_),
    .A2(_1034_),
    .Y(_1037_),
    .B1(_1033_));
 sg13g2_o21ai_1 _4067_ (.B1(_1025_),
    .VDD(VPWR),
    .Y(_1038_),
    .VSS(VGND),
    .A1(_1024_),
    .A2(_1028_));
 sg13g2_xnor2_1 _4068_ (.Y(_1039_),
    .A(net940),
    .B(_1038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4069_ (.Y(_1040_),
    .A(_1030_),
    .B(_1039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4070_ (.Y(_1041_),
    .A(_1037_),
    .B(_1040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4071_ (.B1(net464),
    .VDD(VPWR),
    .Y(_1042_),
    .VSS(VGND),
    .A1(net566),
    .A2(net940));
 sg13g2_a21oi_1 _4072_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net571),
    .A2(_1041_),
    .Y(_0147_),
    .B1(_1042_));
 sg13g2_nand3_1 _4073_ (.B(\mydesign.inputs[1][8] ),
    .C(net460),
    .A(net498),
    .Y(_1043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4074_ (.X(_1044_),
    .A(net544),
    .B(net555),
    .C(\mydesign.inputs[1][12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4075_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\mydesign.inputs[1][20] ),
    .C1(_1044_),
    .B1(net461),
    .A1(\mydesign.inputs[1][16] ),
    .Y(_1045_),
    .A2(net495));
 sg13g2_o21ai_1 _4076_ (.B1(_1043_),
    .VDD(VPWR),
    .Y(_1046_),
    .VSS(VGND),
    .A1(net543),
    .A2(_1045_));
 sg13g2_o21ai_1 _4077_ (.B1(net626),
    .VDD(VPWR),
    .Y(_1047_),
    .VSS(VGND),
    .A1(net489),
    .A2(_1046_));
 sg13g2_a21oi_1 _4078_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2571_),
    .A2(net488),
    .Y(_0148_),
    .B1(_1047_));
 sg13g2_nand3_1 _4079_ (.B(\mydesign.inputs[1][9] ),
    .C(net460),
    .A(net498),
    .Y(_1048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4080_ (.X(_1049_),
    .A(net544),
    .B(net554),
    .C(\mydesign.inputs[1][13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4081_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\mydesign.inputs[1][21] ),
    .C1(_1049_),
    .B1(net461),
    .A1(\mydesign.inputs[1][17] ),
    .Y(_1050_),
    .A2(net495));
 sg13g2_o21ai_1 _4082_ (.B1(_1048_),
    .VDD(VPWR),
    .Y(_1051_),
    .VSS(VGND),
    .A1(net542),
    .A2(_1050_));
 sg13g2_o21ai_1 _4083_ (.B1(net626),
    .VDD(VPWR),
    .Y(_1052_),
    .VSS(VGND),
    .A1(net489),
    .A2(_1051_));
 sg13g2_a21oi_1 _4084_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2570_),
    .A2(net488),
    .Y(_0149_),
    .B1(_1052_));
 sg13g2_nand2_1 _4085_ (.Y(_1053_),
    .A(\mydesign.inputs[1][18] ),
    .B(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4086_ (.Y(_1054_),
    .B1(_0394_),
    .B2(\mydesign.inputs[1][14] ),
    .A2(net461),
    .A1(\mydesign.inputs[1][22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4087_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1053_),
    .A2(_1054_),
    .Y(_1055_),
    .B1(net542));
 sg13g2_a21o_2 _4088_ (.A2(_0639_),
    .A1(net791),
    .B1(_1055_),
    .X(_1056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4089_ (.B1(net626),
    .VDD(VPWR),
    .Y(_1057_),
    .VSS(VGND),
    .A1(net489),
    .A2(_1056_));
 sg13g2_a21oi_1 _4090_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2569_),
    .A2(net489),
    .Y(_0150_),
    .B1(_1057_));
 sg13g2_nand2_1 _4091_ (.Y(_1058_),
    .A(\mydesign.inputs[1][15] ),
    .B(_0394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4092_ (.Y(_1059_),
    .B1(_0390_),
    .B2(\mydesign.inputs[1][23] ),
    .A2(_2595_),
    .A1(\mydesign.inputs[1][19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4093_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1058_),
    .A2(_1059_),
    .Y(_1060_),
    .B1(net542));
 sg13g2_a21o_2 _4094_ (.A2(_0639_),
    .A1(net800),
    .B1(_1060_),
    .X(_1061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4095_ (.B1(net626),
    .VDD(VPWR),
    .Y(_1062_),
    .VSS(VGND),
    .A1(net489),
    .A2(_1061_));
 sg13g2_a21oi_1 _4096_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2568_),
    .A2(net488),
    .Y(_0151_),
    .B1(_1062_));
 sg13g2_o21ai_1 _4097_ (.B1(net624),
    .VDD(VPWR),
    .Y(_1063_),
    .VSS(VGND),
    .A1(net815),
    .A2(net436));
 sg13g2_a21oi_1 _4098_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2578_),
    .A2(net436),
    .Y(_0152_),
    .B1(_1063_));
 sg13g2_o21ai_1 _4099_ (.B1(net624),
    .VDD(VPWR),
    .Y(_1064_),
    .VSS(VGND),
    .A1(net811),
    .A2(net436));
 sg13g2_a21oi_1 _4100_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2577_),
    .A2(net436),
    .Y(_0153_),
    .B1(_1064_));
 sg13g2_o21ai_1 _4101_ (.B1(net624),
    .VDD(VPWR),
    .Y(_1065_),
    .VSS(VGND),
    .A1(\mydesign.pe_weights[46] ),
    .A2(net436));
 sg13g2_a21oi_1 _4102_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2576_),
    .A2(net436),
    .Y(_0154_),
    .B1(_1065_));
 sg13g2_o21ai_1 _4103_ (.B1(net624),
    .VDD(VPWR),
    .Y(_1066_),
    .VSS(VGND),
    .A1(net927),
    .A2(net436));
 sg13g2_a21oi_1 _4104_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2575_),
    .A2(net437),
    .Y(_0155_),
    .B1(_1066_));
 sg13g2_and2_1 _4105_ (.A(net808),
    .B(_1046_),
    .X(_1067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4106_ (.Y(_1068_),
    .A(net561),
    .B(_1067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4107_ (.B(_1068_),
    .A(net1003),
    .X(_1069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4108_ (.A(net462),
    .B(_1069_),
    .Y(_0156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4109_ (.B(\mydesign.pe_weights[61] ),
    .C(_1046_),
    .A(\mydesign.accum[89] ),
    .Y(_1070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4110_ (.A2(_1046_),
    .A1(\mydesign.pe_weights[61] ),
    .B1(\mydesign.accum[89] ),
    .X(_1071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4111_ (.Y(_1072_),
    .A(_1070_),
    .B(_1071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4112_ (.Y(_1073_),
    .A(net808),
    .B(_1051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4113_ (.A(_1072_),
    .B(_1073_),
    .Y(_1074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4114_ (.B(_1073_),
    .A(_1072_),
    .X(_1075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4115_ (.X(_1076_),
    .A(\mydesign.accum[88] ),
    .B(_1067_),
    .C(_1075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4116_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[88] ),
    .A2(_1067_),
    .Y(_1077_),
    .B1(_1075_));
 sg13g2_or2_1 _4117_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1078_),
    .B(_1077_),
    .A(_1076_));
 sg13g2_o21ai_1 _4118_ (.B1(net468),
    .VDD(VPWR),
    .Y(_1079_),
    .VSS(VGND),
    .A1(net561),
    .A2(net896));
 sg13g2_a21oi_1 _4119_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net561),
    .A2(_1078_),
    .Y(_0157_),
    .B1(_1079_));
 sg13g2_nand2_1 _4120_ (.Y(_1080_),
    .A(\mydesign.pe_weights[60] ),
    .B(_1056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4121_ (.X(_1081_),
    .A(\mydesign.accum[90] ),
    .B(\mydesign.pe_weights[62] ),
    .C(_1046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4122_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[62] ),
    .A2(_1046_),
    .Y(_1082_),
    .B1(\mydesign.accum[90] ));
 sg13g2_nand2_1 _4123_ (.Y(_1083_),
    .A(\mydesign.pe_weights[61] ),
    .B(_1051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4124_ (.A(_1081_),
    .B(_1082_),
    .C(_1083_),
    .Y(_1084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4125_ (.B1(_1083_),
    .VDD(VPWR),
    .Y(_1085_),
    .VSS(VGND),
    .A1(_1081_),
    .A2(_1082_));
 sg13g2_nor2b_1 _4126_ (.A(_1084_),
    .B_N(_1085_),
    .Y(_1086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4127_ (.Y(_1087_),
    .B(_1086_),
    .A_N(_1070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4128_ (.Y(_1088_),
    .A(_1070_),
    .B(_1086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4129_ (.Y(_1089_),
    .B(_1088_),
    .A_N(_1080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4130_ (.Y(_1090_),
    .A(_1080_),
    .B(_1088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4131_ (.A(_1074_),
    .B(_1090_),
    .X(_1091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4132_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1092_),
    .B(_1090_),
    .A(_1074_));
 sg13g2_nand2b_1 _4133_ (.Y(_1093_),
    .B(_1092_),
    .A_N(_1091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4134_ (.B(_1093_),
    .A(_1076_),
    .X(_1094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4135_ (.B1(net468),
    .VDD(VPWR),
    .Y(_1095_),
    .VSS(VGND),
    .A1(net560),
    .A2(net964));
 sg13g2_a21oi_1 _4136_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net561),
    .A2(_1094_),
    .Y(_0158_),
    .B1(_1095_));
 sg13g2_a21oi_1 _4137_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1076_),
    .A2(_1092_),
    .Y(_1096_),
    .B1(_1091_));
 sg13g2_nand2_1 _4138_ (.Y(_1097_),
    .A(_1087_),
    .B(_1089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4139_ (.Y(_1098_),
    .A(\mydesign.pe_weights[60] ),
    .B(_1061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4140_ (.VDD(VPWR),
    .Y(_1099_),
    .A(_1098_),
    .VSS(VGND));
 sg13g2_nand2_1 _4141_ (.Y(_1100_),
    .A(\mydesign.pe_weights[61] ),
    .B(_1056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4142_ (.Y(_1101_),
    .A(\mydesign.pe_weights[62] ),
    .B(_1051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4143_ (.X(_1102_),
    .A(\mydesign.accum[91] ),
    .B(\mydesign.pe_weights[63] ),
    .C(_1046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4144_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[63] ),
    .A2(_1046_),
    .Y(_1103_),
    .B1(\mydesign.accum[91] ));
 sg13g2_or3_1 _4145_ (.A(_1101_),
    .B(_1102_),
    .C(_1103_),
    .X(_1104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4146_ (.B1(_1101_),
    .VDD(VPWR),
    .Y(_1105_),
    .VSS(VGND),
    .A1(_1102_),
    .A2(_1103_));
 sg13g2_and3_1 _4147_ (.X(_1106_),
    .A(_1081_),
    .B(_1104_),
    .C(_1105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4148_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1104_),
    .A2(_1105_),
    .Y(_1107_),
    .B1(_1081_));
 sg13g2_or3_1 _4149_ (.A(_1100_),
    .B(_1106_),
    .C(_1107_),
    .X(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4150_ (.B1(_1100_),
    .VDD(VPWR),
    .Y(_1109_),
    .VSS(VGND),
    .A1(_1106_),
    .A2(_1107_));
 sg13g2_nand3_1 _4151_ (.B(_1108_),
    .C(_1109_),
    .A(_1084_),
    .Y(_1110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4152_ (.A2(_1109_),
    .A1(_1108_),
    .B1(_1084_),
    .X(_1111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4153_ (.B(_1110_),
    .C(_1111_),
    .A(_1099_),
    .Y(_1112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4154_ (.A2(_1111_),
    .A1(_1110_),
    .B1(_1099_),
    .X(_1113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4155_ (.X(_1114_),
    .A(_1097_),
    .B(_1112_),
    .C(_1113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4156_ (.B(_1112_),
    .C(_1113_),
    .A(_1097_),
    .Y(_1115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4157_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1112_),
    .A2(_1113_),
    .Y(_1116_),
    .B1(_1097_));
 sg13g2_nor2_1 _4158_ (.A(_1114_),
    .B(_1116_),
    .Y(_1117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4159_ (.Y(_1118_),
    .A(_1096_),
    .B(_1117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4160_ (.B1(net469),
    .VDD(VPWR),
    .Y(_1119_),
    .VSS(VGND),
    .A1(net499),
    .A2(_1118_));
 sg13g2_a21oi_1 _4161_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net500),
    .A2(_2574_),
    .Y(_0159_),
    .B1(_1119_));
 sg13g2_nor2b_1 _4162_ (.A(_1106_),
    .B_N(_1108_),
    .Y(_1120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4163_ (.Y(_1121_),
    .A(\mydesign.pe_weights[61] ),
    .B(_1061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4164_ (.Y(_1122_),
    .B(_1104_),
    .A_N(_1102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4165_ (.Y(_1123_),
    .A(\mydesign.pe_weights[62] ),
    .B(_1056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4166_ (.A(\mydesign.pe_weights[63] ),
    .B(_1051_),
    .X(_1124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4167_ (.Y(_1125_),
    .A(\mydesign.accum[92] ),
    .B(_1124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4168_ (.A(_1123_),
    .B(_1125_),
    .Y(_1126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4169_ (.B(_1125_),
    .A(_1123_),
    .X(_1127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4170_ (.Y(_1128_),
    .A(_1122_),
    .B(_1127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4171_ (.Y(_1129_),
    .A(_1122_),
    .B(_1127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4172_ (.B(_1129_),
    .A(_1121_),
    .X(_1130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4173_ (.Y(_1131_),
    .B(_1130_),
    .A_N(_1120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4174_ (.B(_1130_),
    .A(_1120_),
    .X(_1132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4175_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1110_),
    .A2(_1112_),
    .Y(_1133_),
    .B1(_1132_));
 sg13g2_nand3_1 _4176_ (.B(_1112_),
    .C(_1132_),
    .A(_1110_),
    .Y(_1134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4177_ (.Y(_1135_),
    .B(_1134_),
    .A_N(_1133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4178_ (.B1(_1115_),
    .VDD(VPWR),
    .Y(_1136_),
    .VSS(VGND),
    .A1(_1096_),
    .A2(_1116_));
 sg13g2_xor2_1 _4179_ (.B(_1136_),
    .A(_1135_),
    .X(_1137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4180_ (.B1(net468),
    .VDD(VPWR),
    .Y(_1138_),
    .VSS(VGND),
    .A1(net569),
    .A2(net997));
 sg13g2_a21oi_1 _4181_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net569),
    .A2(_1137_),
    .Y(_0160_),
    .B1(_1138_));
 sg13g2_a21oi_1 _4182_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1134_),
    .A2(_1136_),
    .Y(_1139_),
    .B1(_1133_));
 sg13g2_o21ai_1 _4183_ (.B1(_1128_),
    .VDD(VPWR),
    .Y(_1140_),
    .VSS(VGND),
    .A1(_1121_),
    .A2(_1129_));
 sg13g2_nand2_1 _4184_ (.Y(_1141_),
    .A(\mydesign.pe_weights[62] ),
    .B(_1061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4185_ (.Y(_1142_),
    .A(\mydesign.pe_weights[63] ),
    .B(_1056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4186_ (.Y(_1143_),
    .A(\mydesign.accum[93] ),
    .B(_1142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4187_ (.Y(_1144_),
    .B(_1143_),
    .A_N(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4188_ (.Y(_1145_),
    .A(_1141_),
    .B(_1143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4189_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[92] ),
    .A2(_1124_),
    .Y(_1146_),
    .B1(_1126_));
 sg13g2_nand2b_1 _4190_ (.Y(_1147_),
    .B(_1145_),
    .A_N(_1146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4191_ (.Y(_1148_),
    .A(_1145_),
    .B(_1146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4192_ (.Y(_1149_),
    .A(_1140_),
    .B(_1148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4193_ (.Y(_1150_),
    .A(_1140_),
    .B(_1148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4194_ (.A(_1131_),
    .B(_1150_),
    .X(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4195_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1152_),
    .B(_1150_),
    .A(_1131_));
 sg13g2_nor2b_1 _4196_ (.A(_1151_),
    .B_N(_1152_),
    .Y(_1153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4197_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1154_),
    .B(_1153_),
    .A(_1139_));
 sg13g2_a21oi_1 _4198_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1139_),
    .A2(_1153_),
    .Y(_1155_),
    .B1(net500));
 sg13g2_a221oi_1 _4199_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1155_),
    .C1(net462),
    .B1(_1154_),
    .A1(net500),
    .Y(_0161_),
    .A2(_2573_));
 sg13g2_o21ai_1 _4200_ (.B1(_1144_),
    .VDD(VPWR),
    .Y(_1156_),
    .VSS(VGND),
    .A1(_2573_),
    .A2(_1142_));
 sg13g2_nand2_1 _4201_ (.Y(_1157_),
    .A(\mydesign.pe_weights[63] ),
    .B(_1061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4202_ (.Y(_1158_),
    .A(_2572_),
    .B(_1157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4203_ (.Y(_1159_),
    .B(_1156_),
    .A_N(_1158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4204_ (.B(_1158_),
    .A(_1156_),
    .X(_1160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4205_ (.A(_1147_),
    .B(_1160_),
    .Y(_1161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4206_ (.A(_1149_),
    .B(_1160_),
    .Y(_1162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4207_ (.Y(_1163_),
    .A(_1147_),
    .B(_1149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4208_ (.Y(_1164_),
    .A(_1160_),
    .B(_1163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4209_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1139_),
    .A2(_1152_),
    .Y(_1165_),
    .B1(_1151_));
 sg13g2_xnor2_1 _4210_ (.Y(_1166_),
    .A(_1164_),
    .B(_1165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4211_ (.B1(net471),
    .VDD(VPWR),
    .Y(_1167_),
    .VSS(VGND),
    .A1(net569),
    .A2(net806));
 sg13g2_a21oi_1 _4212_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net569),
    .A2(_1166_),
    .Y(_0162_),
    .B1(_1167_));
 sg13g2_a21oi_1 _4213_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1164_),
    .A2(_1165_),
    .Y(_1168_),
    .B1(_1162_));
 sg13g2_o21ai_1 _4214_ (.B1(_1159_),
    .VDD(VPWR),
    .Y(_1169_),
    .VSS(VGND),
    .A1(_2572_),
    .A2(_1157_));
 sg13g2_xor2_1 _4215_ (.B(_1169_),
    .A(net948),
    .X(_1170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4216_ (.Y(_1171_),
    .A(_1161_),
    .B(_1170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4217_ (.Y(_1172_),
    .A(_1168_),
    .B(_1171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4218_ (.B1(net471),
    .VDD(VPWR),
    .Y(_1173_),
    .VSS(VGND),
    .A1(net569),
    .A2(net948));
 sg13g2_a21oi_1 _4219_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net569),
    .A2(_1172_),
    .Y(_0163_),
    .B1(_1173_));
 sg13g2_o21ai_1 _4220_ (.B1(net631),
    .VDD(VPWR),
    .Y(_1174_),
    .VSS(VGND),
    .A1(net1050),
    .A2(net447));
 sg13g2_a21oi_1 _4221_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2571_),
    .A2(net447),
    .Y(_0164_),
    .B1(_1174_));
 sg13g2_o21ai_1 _4222_ (.B1(net630),
    .VDD(VPWR),
    .Y(_1175_),
    .VSS(VGND),
    .A1(net899),
    .A2(net438));
 sg13g2_a21oi_1 _4223_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2570_),
    .A2(net438),
    .Y(_0165_),
    .B1(_1175_));
 sg13g2_o21ai_1 _4224_ (.B1(net626),
    .VDD(VPWR),
    .Y(_1176_),
    .VSS(VGND),
    .A1(net981),
    .A2(net438));
 sg13g2_a21oi_1 _4225_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2569_),
    .A2(net439),
    .Y(_0166_),
    .B1(_1176_));
 sg13g2_o21ai_1 _4226_ (.B1(net630),
    .VDD(VPWR),
    .Y(_1177_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[43] ),
    .A2(net438));
 sg13g2_a21oi_1 _4227_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2568_),
    .A2(net438),
    .Y(_0167_),
    .B1(_1177_));
 sg13g2_o21ai_1 _4228_ (.B1(net631),
    .VDD(VPWR),
    .Y(_1178_),
    .VSS(VGND),
    .A1(net1013),
    .A2(net447));
 sg13g2_a21oi_1 _4229_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2567_),
    .A2(net447),
    .Y(_0168_),
    .B1(_1178_));
 sg13g2_o21ai_1 _4230_ (.B1(net631),
    .VDD(VPWR),
    .Y(_1179_),
    .VSS(VGND),
    .A1(net856),
    .A2(net448));
 sg13g2_a21oi_1 _4231_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2566_),
    .A2(net448),
    .Y(_0169_),
    .B1(_1179_));
 sg13g2_o21ai_1 _4232_ (.B1(net631),
    .VDD(VPWR),
    .Y(_1180_),
    .VSS(VGND),
    .A1(net813),
    .A2(net448));
 sg13g2_a21oi_1 _4233_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2565_),
    .A2(net448),
    .Y(_0170_),
    .B1(_1180_));
 sg13g2_o21ai_1 _4234_ (.B1(net631),
    .VDD(VPWR),
    .Y(_1181_),
    .VSS(VGND),
    .A1(net533),
    .A2(net448));
 sg13g2_a21oi_1 _4235_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2564_),
    .A2(net448),
    .Y(_0171_),
    .B1(_1181_));
 sg13g2_nor3_1 _4236_ (.A(net502),
    .B(_2567_),
    .C(_2571_),
    .Y(_1182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4237_ (.B1(net479),
    .VDD(VPWR),
    .Y(_1183_),
    .VSS(VGND),
    .A1(net739),
    .A2(_1182_));
 sg13g2_a21oi_1 _4238_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net739),
    .A2(_1182_),
    .Y(_0172_),
    .B1(_1183_));
 sg13g2_and3_2 _4239_ (.X(_1184_),
    .A(\mydesign.accum[81] ),
    .B(\mydesign.pe_weights[57] ),
    .C(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4240_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[57] ),
    .A2(net536),
    .Y(_1185_),
    .B1(\mydesign.accum[81] ));
 sg13g2_nand2_1 _4241_ (.Y(_1186_),
    .A(\mydesign.pe_weights[56] ),
    .B(\mydesign.pe_inputs[45] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4242_ (.A(_1184_),
    .B(_1185_),
    .C(_1186_),
    .Y(_1187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4243_ (.B1(_1186_),
    .VDD(VPWR),
    .Y(_1188_),
    .VSS(VGND),
    .A1(_1184_),
    .A2(_1185_));
 sg13g2_nor2b_1 _4244_ (.A(_1187_),
    .B_N(_1188_),
    .Y(_1189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4245_ (.B(\mydesign.pe_weights[56] ),
    .C(net536),
    .A(net739),
    .Y(_1190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4246_ (.B(\mydesign.pe_weights[56] ),
    .C(net536),
    .A(net739),
    .Y(_1191_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1189_));
 sg13g2_xor2_1 _4247_ (.B(_1190_),
    .A(_1189_),
    .X(_1192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4248_ (.B1(net471),
    .VDD(VPWR),
    .Y(_1193_),
    .VSS(VGND),
    .A1(net570),
    .A2(net983));
 sg13g2_a21oi_1 _4249_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net570),
    .A2(_1192_),
    .Y(_0173_),
    .B1(_1193_));
 sg13g2_nand2_1 _4250_ (.Y(_1194_),
    .A(\mydesign.pe_weights[56] ),
    .B(\mydesign.pe_inputs[46] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4251_ (.Y(_1195_),
    .A(\mydesign.pe_weights[57] ),
    .B(\mydesign.pe_inputs[45] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4252_ (.B(\mydesign.pe_weights[58] ),
    .C(net536),
    .A(\mydesign.accum[82] ),
    .Y(_1196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4253_ (.A2(net536),
    .A1(\mydesign.pe_weights[58] ),
    .B1(\mydesign.accum[82] ),
    .X(_1197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4254_ (.Y(_1198_),
    .A(_1196_),
    .B(_1197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4255_ (.A(_1195_),
    .B(_1198_),
    .Y(_1199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4256_ (.B(_1198_),
    .A(_1195_),
    .X(_1200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4257_ (.Y(_1201_),
    .A(_1184_),
    .B(_1200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4258_ (.A(_1184_),
    .B(_1200_),
    .Y(_1202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4259_ (.B(_1200_),
    .A(_1184_),
    .X(_1203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4260_ (.Y(_1204_),
    .A(_1194_),
    .B(_1203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4261_ (.Y(_1205_),
    .A(_1187_),
    .B(_1204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4262_ (.Y(_1206_),
    .A(_1187_),
    .B(_1204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4263_ (.Y(_1207_),
    .A(_1191_),
    .B(_1206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4264_ (.B1(net472),
    .VDD(VPWR),
    .Y(_1208_),
    .VSS(VGND),
    .A1(net570),
    .A2(net961));
 sg13g2_a21oi_1 _4265_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net570),
    .A2(_1207_),
    .Y(_0174_),
    .B1(_1208_));
 sg13g2_o21ai_1 _4266_ (.B1(_1205_),
    .VDD(VPWR),
    .Y(_1209_),
    .VSS(VGND),
    .A1(_1191_),
    .A2(_1206_));
 sg13g2_o21ai_1 _4267_ (.B1(_1201_),
    .VDD(VPWR),
    .Y(_1210_),
    .VSS(VGND),
    .A1(_1194_),
    .A2(_1202_));
 sg13g2_nand2_1 _4268_ (.Y(_1211_),
    .A(\mydesign.pe_weights[56] ),
    .B(\mydesign.pe_inputs[47] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4269_ (.Y(_1212_),
    .A(\mydesign.pe_weights[57] ),
    .B(\mydesign.pe_inputs[46] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4270_ (.Y(_1213_),
    .A(\mydesign.pe_weights[58] ),
    .B(\mydesign.pe_inputs[45] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4271_ (.B(net539),
    .C(net536),
    .A(\mydesign.accum[83] ),
    .Y(_1214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4272_ (.A2(\mydesign.pe_inputs[44] ),
    .A1(net539),
    .B1(\mydesign.accum[83] ),
    .X(_1215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4273_ (.Y(_1216_),
    .A(_1214_),
    .B(_1215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4274_ (.B(_1216_),
    .A(_1213_),
    .X(_1217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4275_ (.A(_1196_),
    .B_N(_1217_),
    .Y(_1218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4276_ (.B(_1217_),
    .A(_1196_),
    .X(_1219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4277_ (.A(_1212_),
    .B(_1219_),
    .Y(_1220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4278_ (.B(_1219_),
    .A(_1212_),
    .X(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4279_ (.Y(_1222_),
    .A(_1199_),
    .B(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4280_ (.Y(_1223_),
    .A(_1199_),
    .B(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4281_ (.B(_1223_),
    .A(_1211_),
    .X(_1224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4282_ (.A(_1210_),
    .B(_1224_),
    .X(_1225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4283_ (.Y(_1226_),
    .A(_1210_),
    .B(_1224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4284_ (.A(_1226_),
    .B_N(_1209_),
    .Y(_1227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4285_ (.B(_1226_),
    .A(_1209_),
    .X(_1228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4286_ (.B1(net471),
    .VDD(VPWR),
    .Y(_1229_),
    .VSS(VGND),
    .A1(net579),
    .A2(net911));
 sg13g2_a21oi_1 _4287_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net579),
    .A2(_1228_),
    .Y(_0175_),
    .B1(_1229_));
 sg13g2_nand2_1 _4288_ (.Y(_1230_),
    .A(\mydesign.pe_weights[57] ),
    .B(\mydesign.pe_inputs[47] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4289_ (.B1(_1214_),
    .VDD(VPWR),
    .Y(_1231_),
    .VSS(VGND),
    .A1(_1213_),
    .A2(_1216_));
 sg13g2_nand2_1 _4290_ (.Y(_1232_),
    .A(\mydesign.pe_weights[58] ),
    .B(\mydesign.pe_inputs[46] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4291_ (.B(net539),
    .C(\mydesign.pe_inputs[45] ),
    .A(\mydesign.accum[84] ),
    .Y(_1233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4292_ (.A2(\mydesign.pe_inputs[45] ),
    .A1(net539),
    .B1(\mydesign.accum[84] ),
    .X(_1234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4293_ (.Y(_1235_),
    .A(_1233_),
    .B(_1234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4294_ (.B(_1235_),
    .A(_1232_),
    .X(_1236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4295_ (.Y(_1237_),
    .A(_1231_),
    .B(_1236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4296_ (.Y(_1238_),
    .A(_1231_),
    .B(_1236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4297_ (.B(_1238_),
    .A(_1230_),
    .X(_1239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4298_ (.B1(_1239_),
    .VDD(VPWR),
    .Y(_1240_),
    .VSS(VGND),
    .A1(_1218_),
    .A2(_1220_));
 sg13g2_or3_1 _4299_ (.A(_1218_),
    .B(_1220_),
    .C(_1239_),
    .X(_1241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4300_ (.A(_1240_),
    .B(_1241_),
    .X(_1242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4301_ (.B1(_1222_),
    .VDD(VPWR),
    .Y(_1243_),
    .VSS(VGND),
    .A1(_1211_),
    .A2(_1223_));
 sg13g2_nand2_1 _4302_ (.Y(_1244_),
    .A(_1242_),
    .B(_1243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4303_ (.B(_1243_),
    .A(_1242_),
    .X(_1245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4304_ (.A(_1225_),
    .B(_1227_),
    .C(_1245_),
    .Y(_1246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4305_ (.B1(_1245_),
    .VDD(VPWR),
    .Y(_1247_),
    .VSS(VGND),
    .A1(_1225_),
    .A2(_1227_));
 sg13g2_nand2b_1 _4306_ (.Y(_1248_),
    .B(_1247_),
    .A_N(_1246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4307_ (.B1(net471),
    .VDD(VPWR),
    .Y(_1249_),
    .VSS(VGND),
    .A1(net579),
    .A2(net933));
 sg13g2_a21oi_1 _4308_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net579),
    .A2(_1248_),
    .Y(_0176_),
    .B1(_1249_));
 sg13g2_nand2_1 _4309_ (.Y(_1250_),
    .A(\mydesign.pe_weights[58] ),
    .B(\mydesign.pe_inputs[47] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4310_ (.X(_1251_),
    .A(\mydesign.accum[85] ),
    .B(net539),
    .C(\mydesign.pe_inputs[46] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4311_ (.B(\mydesign.pe_weights[59] ),
    .C(\mydesign.pe_inputs[46] ),
    .A(\mydesign.accum[85] ),
    .Y(_1252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4312_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[59] ),
    .A2(\mydesign.pe_inputs[46] ),
    .Y(_1253_),
    .B1(\mydesign.accum[85] ));
 sg13g2_nor2_1 _4313_ (.A(_1251_),
    .B(_1253_),
    .Y(_1254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4314_ (.Y(_1255_),
    .A(_1250_),
    .B(_1254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4315_ (.B1(_1233_),
    .VDD(VPWR),
    .Y(_1256_),
    .VSS(VGND),
    .A1(_1232_),
    .A2(_1235_));
 sg13g2_xor2_1 _4316_ (.B(_1256_),
    .A(_1255_),
    .X(_1257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4317_ (.B1(_1237_),
    .VDD(VPWR),
    .Y(_1258_),
    .VSS(VGND),
    .A1(_1230_),
    .A2(_1238_));
 sg13g2_nand2_1 _4318_ (.Y(_1259_),
    .A(_1257_),
    .B(_1258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4319_ (.B(_1258_),
    .A(_1257_),
    .X(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4320_ (.A(_1240_),
    .B_N(_1260_),
    .Y(_1261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4321_ (.B(_1260_),
    .A(_1240_),
    .X(_1262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4322_ (.X(_1263_),
    .A(_1244_),
    .B(_1247_),
    .C(_1262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4323_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1244_),
    .A2(_1247_),
    .Y(_1264_),
    .B1(_1262_));
 sg13g2_o21ai_1 _4324_ (.B1(net579),
    .VDD(VPWR),
    .Y(_1265_),
    .VSS(VGND),
    .A1(_1263_),
    .A2(_1264_));
 sg13g2_o21ai_1 _4325_ (.B1(net479),
    .VDD(VPWR),
    .Y(_1266_),
    .VSS(VGND),
    .A1(net580),
    .A2(net951));
 sg13g2_nor2b_1 _4326_ (.A(_1266_),
    .B_N(_1265_),
    .Y(_0177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4327_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net539),
    .A2(\mydesign.pe_inputs[47] ),
    .Y(_1267_),
    .B1(\mydesign.accum[86] ));
 sg13g2_nand3_1 _4328_ (.B(net539),
    .C(\mydesign.pe_inputs[47] ),
    .A(\mydesign.accum[86] ),
    .Y(_1268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4329_ (.Y(_1269_),
    .B(_1268_),
    .A_N(_1267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4330_ (.B1(_1252_),
    .VDD(VPWR),
    .Y(_1270_),
    .VSS(VGND),
    .A1(_1250_),
    .A2(_1253_));
 sg13g2_inv_1 _4331_ (.VDD(VPWR),
    .Y(_1271_),
    .A(_1270_),
    .VSS(VGND));
 sg13g2_xnor2_1 _4332_ (.Y(_1272_),
    .A(_1269_),
    .B(_1270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4333_ (.B(_1256_),
    .C(_1272_),
    .A(_1255_),
    .Y(_1273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4334_ (.A2(_1256_),
    .A1(_1255_),
    .B1(_1272_),
    .X(_1274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4335_ (.A(_1273_),
    .B(_1274_),
    .X(_1275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4336_ (.B(_1258_),
    .C(_1275_),
    .A(_1257_),
    .Y(_1276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4337_ (.Y(_1277_),
    .A(_1259_),
    .B(_1275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4338_ (.A(_1261_),
    .B(_1264_),
    .C(_1277_),
    .Y(_1278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4339_ (.B1(_1277_),
    .VDD(VPWR),
    .Y(_1279_),
    .VSS(VGND),
    .A1(_1261_),
    .A2(_1264_));
 sg13g2_nand2b_1 _4340_ (.Y(_1280_),
    .B(_1279_),
    .A_N(_1278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4341_ (.B1(net472),
    .VDD(VPWR),
    .Y(_1281_),
    .VSS(VGND),
    .A1(net579),
    .A2(net895));
 sg13g2_a21oi_1 _4342_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net579),
    .A2(_1280_),
    .Y(_0178_),
    .B1(_1281_));
 sg13g2_nand2_1 _4343_ (.Y(_1282_),
    .A(_1276_),
    .B(_1279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4344_ (.B1(_1268_),
    .VDD(VPWR),
    .Y(_1283_),
    .VSS(VGND),
    .A1(_1267_),
    .A2(_1271_));
 sg13g2_xnor2_1 _4345_ (.Y(_1284_),
    .A(net865),
    .B(_1283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4346_ (.Y(_1285_),
    .A(_1273_),
    .B(_1284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4347_ (.B(_1285_),
    .A(_1282_),
    .X(_1286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4348_ (.B1(net479),
    .VDD(VPWR),
    .Y(_1287_),
    .VSS(VGND),
    .A1(net579),
    .A2(net865));
 sg13g2_a21oi_1 _4349_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net580),
    .A2(_1286_),
    .Y(_0179_),
    .B1(_1287_));
 sg13g2_o21ai_1 _4350_ (.B1(net629),
    .VDD(VPWR),
    .Y(_1288_),
    .VSS(VGND),
    .A1(net532),
    .A2(net440));
 sg13g2_a21oi_1 _4351_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2563_),
    .A2(net440),
    .Y(_0180_),
    .B1(_1288_));
 sg13g2_o21ai_1 _4352_ (.B1(net628),
    .VDD(VPWR),
    .Y(_1289_),
    .VSS(VGND),
    .A1(net966),
    .A2(net434));
 sg13g2_a21oi_1 _4353_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2562_),
    .A2(net433),
    .Y(_0181_),
    .B1(_1289_));
 sg13g2_o21ai_1 _4354_ (.B1(net628),
    .VDD(VPWR),
    .Y(_1290_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[38] ),
    .A2(net434));
 sg13g2_a21oi_1 _4355_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2561_),
    .A2(net434),
    .Y(_0182_),
    .B1(_1290_));
 sg13g2_o21ai_1 _4356_ (.B1(net629),
    .VDD(VPWR),
    .Y(_1291_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[39] ),
    .A2(net434));
 sg13g2_a21oi_1 _4357_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2560_),
    .A2(net434),
    .Y(_0183_),
    .B1(_1291_));
 sg13g2_o21ai_1 _4358_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1292_),
    .VSS(VGND),
    .A1(net943),
    .A2(net446));
 sg13g2_a21oi_1 _4359_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2559_),
    .A2(net446),
    .Y(_0184_),
    .B1(_1292_));
 sg13g2_o21ai_1 _4360_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1293_),
    .VSS(VGND),
    .A1(net862),
    .A2(net441));
 sg13g2_a21oi_1 _4361_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2558_),
    .A2(net441),
    .Y(_0185_),
    .B1(_1293_));
 sg13g2_o21ai_1 _4362_ (.B1(net636),
    .VDD(VPWR),
    .Y(_1294_),
    .VSS(VGND),
    .A1(net830),
    .A2(net441));
 sg13g2_a21oi_1 _4363_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2557_),
    .A2(net441),
    .Y(_0186_),
    .B1(_1294_));
 sg13g2_o21ai_1 _4364_ (.B1(net637),
    .VDD(VPWR),
    .Y(_1295_),
    .VSS(VGND),
    .A1(net538),
    .A2(net493));
 sg13g2_a21oi_1 _4365_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2533_),
    .A2(net493),
    .Y(_0187_),
    .B1(_1295_));
 sg13g2_nor3_1 _4366_ (.A(net501),
    .B(_2559_),
    .C(_2563_),
    .Y(_1296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4367_ (.B1(net473),
    .VDD(VPWR),
    .Y(_1297_),
    .VSS(VGND),
    .A1(net684),
    .A2(_1296_));
 sg13g2_a21oi_1 _4368_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net684),
    .A2(_1296_),
    .Y(_0188_),
    .B1(_1297_));
 sg13g2_and3_2 _4369_ (.X(_1298_),
    .A(\mydesign.accum[73] ),
    .B(\mydesign.pe_weights[53] ),
    .C(net534),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4370_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[53] ),
    .A2(net534),
    .Y(_1299_),
    .B1(\mydesign.accum[73] ));
 sg13g2_nand2_1 _4371_ (.Y(_1300_),
    .A(\mydesign.pe_weights[52] ),
    .B(\mydesign.pe_inputs[41] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4372_ (.A(_1298_),
    .B(_1299_),
    .C(_1300_),
    .Y(_1301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4373_ (.B1(_1300_),
    .VDD(VPWR),
    .Y(_1302_),
    .VSS(VGND),
    .A1(_1298_),
    .A2(_1299_));
 sg13g2_nor2b_1 _4374_ (.A(_1301_),
    .B_N(_1302_),
    .Y(_1303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4375_ (.B(\mydesign.pe_weights[52] ),
    .C(net534),
    .A(net684),
    .Y(_1304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4376_ (.B(\mydesign.pe_weights[52] ),
    .C(net534),
    .A(net684),
    .Y(_1305_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1303_));
 sg13g2_xor2_1 _4377_ (.B(_1304_),
    .A(_1303_),
    .X(_1306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4378_ (.B1(net478),
    .VDD(VPWR),
    .Y(_1307_),
    .VSS(VGND),
    .A1(net573),
    .A2(net875));
 sg13g2_a21oi_1 _4379_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net573),
    .A2(_1306_),
    .Y(_0189_),
    .B1(_1307_));
 sg13g2_nand2_1 _4380_ (.Y(_1308_),
    .A(\mydesign.pe_weights[52] ),
    .B(\mydesign.pe_inputs[42] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4381_ (.Y(_1309_),
    .A(\mydesign.pe_weights[53] ),
    .B(\mydesign.pe_inputs[41] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4382_ (.B(\mydesign.pe_weights[54] ),
    .C(net534),
    .A(\mydesign.accum[74] ),
    .Y(_1310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4383_ (.A2(net534),
    .A1(\mydesign.pe_weights[54] ),
    .B1(\mydesign.accum[74] ),
    .X(_1311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4384_ (.Y(_1312_),
    .A(_1310_),
    .B(_1311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4385_ (.A(_1309_),
    .B(_1312_),
    .Y(_1313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4386_ (.B(_1312_),
    .A(_1309_),
    .X(_1314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4387_ (.Y(_1315_),
    .A(_1298_),
    .B(_1314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4388_ (.A(_1298_),
    .B(_1314_),
    .Y(_1316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4389_ (.B(_1314_),
    .A(_1298_),
    .X(_1317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4390_ (.Y(_1318_),
    .A(_1308_),
    .B(_1317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4391_ (.Y(_1319_),
    .A(_1301_),
    .B(_1318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4392_ (.Y(_1320_),
    .A(_1301_),
    .B(_1318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4393_ (.Y(_1321_),
    .A(_1305_),
    .B(_1320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4394_ (.B1(net474),
    .VDD(VPWR),
    .Y(_1322_),
    .VSS(VGND),
    .A1(net575),
    .A2(net882));
 sg13g2_a21oi_1 _4395_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net575),
    .A2(_1321_),
    .Y(_0190_),
    .B1(_1322_));
 sg13g2_o21ai_1 _4396_ (.B1(_1319_),
    .VDD(VPWR),
    .Y(_1323_),
    .VSS(VGND),
    .A1(_1305_),
    .A2(_1320_));
 sg13g2_o21ai_1 _4397_ (.B1(_1315_),
    .VDD(VPWR),
    .Y(_1324_),
    .VSS(VGND),
    .A1(_1308_),
    .A2(_1316_));
 sg13g2_nand2_1 _4398_ (.Y(_1325_),
    .A(\mydesign.pe_weights[52] ),
    .B(\mydesign.pe_inputs[43] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4399_ (.Y(_1326_),
    .A(\mydesign.pe_weights[53] ),
    .B(\mydesign.pe_inputs[42] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4400_ (.Y(_1327_),
    .A(\mydesign.pe_weights[54] ),
    .B(\mydesign.pe_inputs[41] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4401_ (.B(net538),
    .C(\mydesign.pe_inputs[40] ),
    .A(\mydesign.accum[75] ),
    .Y(_1328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4402_ (.A2(net534),
    .A1(net538),
    .B1(\mydesign.accum[75] ),
    .X(_1329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4403_ (.Y(_1330_),
    .A(_1328_),
    .B(_1329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4404_ (.B(_1330_),
    .A(_1327_),
    .X(_1331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4405_ (.A(_1310_),
    .B_N(_1331_),
    .Y(_1332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4406_ (.B(_1331_),
    .A(_1310_),
    .X(_1333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4407_ (.A(_1326_),
    .B(_1333_),
    .Y(_1334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4408_ (.B(_1333_),
    .A(_1326_),
    .X(_1335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4409_ (.Y(_1336_),
    .A(_1313_),
    .B(_1335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4410_ (.Y(_1337_),
    .A(_1313_),
    .B(_1335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4411_ (.B(_1337_),
    .A(_1325_),
    .X(_1338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4412_ (.A(_1324_),
    .B(_1338_),
    .X(_1339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4413_ (.Y(_1340_),
    .A(_1324_),
    .B(_1338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4414_ (.A(_1340_),
    .B_N(_1323_),
    .Y(_1341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4415_ (.B(_1340_),
    .A(_1323_),
    .X(_1342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4416_ (.B1(net474),
    .VDD(VPWR),
    .Y(_1343_),
    .VSS(VGND),
    .A1(net575),
    .A2(net868));
 sg13g2_a21oi_1 _4417_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net576),
    .A2(_1342_),
    .Y(_0191_),
    .B1(_1343_));
 sg13g2_nand2_1 _4418_ (.Y(_1344_),
    .A(\mydesign.pe_weights[53] ),
    .B(\mydesign.pe_inputs[43] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4419_ (.B1(_1328_),
    .VDD(VPWR),
    .Y(_1345_),
    .VSS(VGND),
    .A1(_1327_),
    .A2(_1330_));
 sg13g2_nand2_1 _4420_ (.Y(_1346_),
    .A(\mydesign.pe_weights[54] ),
    .B(\mydesign.pe_inputs[42] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4421_ (.B(net538),
    .C(\mydesign.pe_inputs[41] ),
    .A(\mydesign.accum[76] ),
    .Y(_1347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4422_ (.A2(\mydesign.pe_inputs[41] ),
    .A1(net538),
    .B1(\mydesign.accum[76] ),
    .X(_1348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4423_ (.Y(_1349_),
    .A(_1347_),
    .B(_1348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4424_ (.B(_1349_),
    .A(_1346_),
    .X(_1350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4425_ (.Y(_1351_),
    .A(_1345_),
    .B(_1350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4426_ (.Y(_1352_),
    .A(_1345_),
    .B(_1350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4427_ (.B(_1352_),
    .A(_1344_),
    .X(_1353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4428_ (.B1(_1353_),
    .VDD(VPWR),
    .Y(_1354_),
    .VSS(VGND),
    .A1(_1332_),
    .A2(_1334_));
 sg13g2_or3_1 _4429_ (.A(_1332_),
    .B(_1334_),
    .C(_1353_),
    .X(_1355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4430_ (.A(_1354_),
    .B(_1355_),
    .X(_1356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4431_ (.B1(_1336_),
    .VDD(VPWR),
    .Y(_1357_),
    .VSS(VGND),
    .A1(_1325_),
    .A2(_1337_));
 sg13g2_nand2_1 _4432_ (.Y(_1358_),
    .A(_1356_),
    .B(_1357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4433_ (.B(_1357_),
    .A(_1356_),
    .X(_1359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4434_ (.A(_1339_),
    .B(_1341_),
    .C(_1359_),
    .X(_1360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4435_ (.B1(_1359_),
    .VDD(VPWR),
    .Y(_1361_),
    .VSS(VGND),
    .A1(_1339_),
    .A2(_1341_));
 sg13g2_a21oi_1 _4436_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1360_),
    .A2(_1361_),
    .Y(_1362_),
    .B1(net501));
 sg13g2_o21ai_1 _4437_ (.B1(net474),
    .VDD(VPWR),
    .Y(_1363_),
    .VSS(VGND),
    .A1(net573),
    .A2(net886));
 sg13g2_nor2_1 _4438_ (.A(_1362_),
    .B(_1363_),
    .Y(_0192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4439_ (.Y(_1364_),
    .A(\mydesign.pe_weights[54] ),
    .B(\mydesign.pe_inputs[43] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4440_ (.B(\mydesign.pe_weights[55] ),
    .C(\mydesign.pe_inputs[42] ),
    .A(\mydesign.accum[77] ),
    .Y(_1365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4441_ (.A2(\mydesign.pe_inputs[42] ),
    .A1(\mydesign.pe_weights[55] ),
    .B1(\mydesign.accum[77] ),
    .X(_1366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4442_ (.Y(_1367_),
    .A(_1365_),
    .B(_1366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4443_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1368_),
    .B(_1367_),
    .A(_1364_));
 sg13g2_xor2_1 _4444_ (.B(_1367_),
    .A(_1364_),
    .X(_1369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4445_ (.B1(_1347_),
    .VDD(VPWR),
    .Y(_1370_),
    .VSS(VGND),
    .A1(_1346_),
    .A2(_1349_));
 sg13g2_and2_1 _4446_ (.A(_1369_),
    .B(_1370_),
    .X(_1371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4447_ (.B(_1370_),
    .A(_1369_),
    .X(_1372_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4448_ (.B1(_1351_),
    .VDD(VPWR),
    .Y(_1373_),
    .VSS(VGND),
    .A1(_1344_),
    .A2(_1352_));
 sg13g2_nand2_1 _4449_ (.Y(_1374_),
    .A(_1372_),
    .B(_1373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4450_ (.B(_1373_),
    .A(_1372_),
    .X(_1375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4451_ (.A(_1354_),
    .B_N(_1375_),
    .Y(_1376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4452_ (.B(_1375_),
    .A(_1354_),
    .X(_1377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4453_ (.X(_1378_),
    .A(_1358_),
    .B(_1361_),
    .C(_1377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4454_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1358_),
    .A2(_1361_),
    .Y(_1379_),
    .B1(_1377_));
 sg13g2_o21ai_1 _4455_ (.B1(net576),
    .VDD(VPWR),
    .Y(_1380_),
    .VSS(VGND),
    .A1(_1378_),
    .A2(_1379_));
 sg13g2_o21ai_1 _4456_ (.B1(_1380_),
    .VDD(VPWR),
    .Y(_1381_),
    .VSS(VGND),
    .A1(net583),
    .A2(net905));
 sg13g2_nor2_1 _4457_ (.A(net463),
    .B(_1381_),
    .Y(_0193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4458_ (.B(net538),
    .C(\mydesign.pe_inputs[43] ),
    .A(\mydesign.accum[78] ),
    .Y(_1382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4459_ (.A2(\mydesign.pe_inputs[43] ),
    .A1(net538),
    .B1(\mydesign.accum[78] ),
    .X(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4460_ (.Y(_1384_),
    .A(_1382_),
    .B(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4461_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1365_),
    .A2(_1368_),
    .Y(_1385_),
    .B1(_1384_));
 sg13g2_nand3_1 _4462_ (.B(_1368_),
    .C(_1384_),
    .A(_1365_),
    .Y(_1386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4463_ (.Y(_1387_),
    .B(_1386_),
    .A_N(_1385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4464_ (.Y(_1388_),
    .B(_1374_),
    .A_N(_1371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4465_ (.Y(_1389_),
    .A(_1387_),
    .B(_1388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4466_ (.A(_1376_),
    .B(_1379_),
    .C(_1389_),
    .X(_1390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4467_ (.B1(_1389_),
    .VDD(VPWR),
    .Y(_1391_),
    .VSS(VGND),
    .A1(_1376_),
    .A2(_1379_));
 sg13g2_a21oi_1 _4468_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1390_),
    .A2(_1391_),
    .Y(_1392_),
    .B1(net502));
 sg13g2_o21ai_1 _4469_ (.B1(net480),
    .VDD(VPWR),
    .Y(_1393_),
    .VSS(VGND),
    .A1(net583),
    .A2(net909));
 sg13g2_nor2_1 _4470_ (.A(_1392_),
    .B(_1393_),
    .Y(_0194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4471_ (.B1(_1391_),
    .VDD(VPWR),
    .Y(_1394_),
    .VSS(VGND),
    .A1(_1374_),
    .A2(_1387_));
 sg13g2_a21oi_1 _4472_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1371_),
    .A2(_1386_),
    .Y(_1395_),
    .B1(_1385_));
 sg13g2_xnor2_1 _4473_ (.Y(_1396_),
    .A(net977),
    .B(_1382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4474_ (.Y(_1397_),
    .A(_1395_),
    .B(_1396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4475_ (.Y(_1398_),
    .A(_1394_),
    .B(_1397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4476_ (.B1(net480),
    .VDD(VPWR),
    .Y(_1399_),
    .VSS(VGND),
    .A1(net581),
    .A2(net977));
 sg13g2_a21oi_1 _4477_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net581),
    .A2(_1398_),
    .Y(_0195_),
    .B1(_1399_));
 sg13g2_nand2b_1 _4478_ (.Y(_1400_),
    .B(_2619_),
    .A_N(_2607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4479_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1401_),
    .B(_1400_),
    .A(_2618_));
 sg13g2_and2_1 _4480_ (.A(net618),
    .B(_1401_),
    .X(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4481_ (.Y(_1403_),
    .A(net646),
    .B(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4482_ (.B1(_1403_),
    .VDD(VPWR),
    .Y(_0196_),
    .VSS(VGND),
    .A1(net603),
    .A2(_1401_));
 sg13g2_nand2_1 _4483_ (.Y(_1404_),
    .A(net644),
    .B(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4484_ (.B1(_1404_),
    .VDD(VPWR),
    .Y(_0197_),
    .VSS(VGND),
    .A1(net601),
    .A2(_1401_));
 sg13g2_nand2_1 _4485_ (.Y(_1405_),
    .A(net422),
    .B(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4486_ (.B1(_1405_),
    .VDD(VPWR),
    .Y(_0198_),
    .VSS(VGND),
    .A1(net599),
    .A2(_1401_));
 sg13g2_nand2_1 _4487_ (.Y(_1406_),
    .A(net666),
    .B(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4488_ (.B1(_1406_),
    .VDD(VPWR),
    .Y(_0199_),
    .VSS(VGND),
    .A1(net597),
    .A2(_1401_));
 sg13g2_o21ai_1 _4489_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1407_),
    .VSS(VGND),
    .A1(\mydesign.pe_weights[48] ),
    .A2(net491));
 sg13g2_a21oi_1 _4490_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2532_),
    .A2(net493),
    .Y(_0200_),
    .B1(_1407_));
 sg13g2_o21ai_1 _4491_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1408_),
    .VSS(VGND),
    .A1(net828),
    .A2(net440));
 sg13g2_a21oi_1 _4492_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2555_),
    .A2(net441),
    .Y(_0201_),
    .B1(_1408_));
 sg13g2_o21ai_1 _4493_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1409_),
    .VSS(VGND),
    .A1(net530),
    .A2(net440));
 sg13g2_a21oi_1 _4494_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2554_),
    .A2(net440),
    .Y(_0202_),
    .B1(_1409_));
 sg13g2_o21ai_1 _4495_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1410_),
    .VSS(VGND),
    .A1(net816),
    .A2(net440));
 sg13g2_a21oi_1 _4496_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2553_),
    .A2(net441),
    .Y(_0203_),
    .B1(_1410_));
 sg13g2_and3_1 _4497_ (.X(_1411_),
    .A(net575),
    .B(\mydesign.pe_weights[48] ),
    .C(net532),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4498_ (.B1(net473),
    .VDD(VPWR),
    .Y(_1412_),
    .VSS(VGND),
    .A1(net690),
    .A2(_1411_));
 sg13g2_a21oi_1 _4499_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net690),
    .A2(_1411_),
    .Y(_0204_),
    .B1(_1412_));
 sg13g2_and3_2 _4500_ (.X(_1413_),
    .A(\mydesign.accum[65] ),
    .B(\mydesign.pe_weights[49] ),
    .C(net532),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4501_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[49] ),
    .A2(net532),
    .Y(_1414_),
    .B1(\mydesign.accum[65] ));
 sg13g2_nand2_1 _4502_ (.Y(_1415_),
    .A(\mydesign.pe_weights[48] ),
    .B(\mydesign.pe_inputs[37] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4503_ (.A(_1413_),
    .B(_1414_),
    .C(_1415_),
    .Y(_1416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4504_ (.B1(_1415_),
    .VDD(VPWR),
    .Y(_1417_),
    .VSS(VGND),
    .A1(_1413_),
    .A2(_1414_));
 sg13g2_nor2b_1 _4505_ (.A(_1416_),
    .B_N(_1417_),
    .Y(_1418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4506_ (.B(\mydesign.pe_weights[48] ),
    .C(\mydesign.pe_inputs[36] ),
    .A(net690),
    .Y(_1419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4507_ (.B(\mydesign.pe_weights[48] ),
    .C(\mydesign.pe_inputs[36] ),
    .A(net690),
    .Y(_1420_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1418_));
 sg13g2_xor2_1 _4508_ (.B(_1419_),
    .A(_1418_),
    .X(_1421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4509_ (.B1(net473),
    .VDD(VPWR),
    .Y(_1422_),
    .VSS(VGND),
    .A1(net574),
    .A2(net907));
 sg13g2_a21oi_1 _4510_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net574),
    .A2(_1421_),
    .Y(_0205_),
    .B1(_1422_));
 sg13g2_nand2_1 _4511_ (.Y(_1423_),
    .A(\mydesign.pe_weights[48] ),
    .B(\mydesign.pe_inputs[38] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4512_ (.Y(_1424_),
    .A(\mydesign.pe_weights[49] ),
    .B(\mydesign.pe_inputs[37] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4513_ (.B(\mydesign.pe_weights[50] ),
    .C(net532),
    .A(\mydesign.accum[66] ),
    .Y(_1425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4514_ (.A2(net532),
    .A1(\mydesign.pe_weights[50] ),
    .B1(\mydesign.accum[66] ),
    .X(_1426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4515_ (.Y(_1427_),
    .A(_1425_),
    .B(_1426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4516_ (.A(_1424_),
    .B(_1427_),
    .Y(_1428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4517_ (.B(_1427_),
    .A(_1424_),
    .X(_1429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4518_ (.Y(_1430_),
    .A(_1413_),
    .B(_1429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4519_ (.A(_1413_),
    .B(_1429_),
    .Y(_1431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4520_ (.B(_1429_),
    .A(_1413_),
    .X(_1432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4521_ (.Y(_1433_),
    .A(_1423_),
    .B(_1432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4522_ (.Y(_1434_),
    .A(_1416_),
    .B(_1433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4523_ (.Y(_1435_),
    .A(_1416_),
    .B(_1433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4524_ (.Y(_1436_),
    .A(_1420_),
    .B(_1435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4525_ (.B1(net464),
    .VDD(VPWR),
    .Y(_1437_),
    .VSS(VGND),
    .A1(net566),
    .A2(net873));
 sg13g2_a21oi_1 _4526_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net566),
    .A2(_1436_),
    .Y(_0206_),
    .B1(_1437_));
 sg13g2_o21ai_1 _4527_ (.B1(_1434_),
    .VDD(VPWR),
    .Y(_1438_),
    .VSS(VGND),
    .A1(_1420_),
    .A2(_1435_));
 sg13g2_o21ai_1 _4528_ (.B1(_1430_),
    .VDD(VPWR),
    .Y(_1439_),
    .VSS(VGND),
    .A1(_1423_),
    .A2(_1431_));
 sg13g2_nand2_1 _4529_ (.Y(_1440_),
    .A(\mydesign.pe_weights[48] ),
    .B(\mydesign.pe_inputs[39] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4530_ (.Y(_1441_),
    .A(\mydesign.pe_weights[49] ),
    .B(\mydesign.pe_inputs[38] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4531_ (.Y(_1442_),
    .A(\mydesign.pe_weights[50] ),
    .B(\mydesign.pe_inputs[37] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4532_ (.B(net537),
    .C(net532),
    .A(\mydesign.accum[67] ),
    .Y(_1443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4533_ (.A2(net532),
    .A1(net537),
    .B1(\mydesign.accum[67] ),
    .X(_1444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4534_ (.Y(_1445_),
    .A(_1443_),
    .B(_1444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4535_ (.B(_1445_),
    .A(_1442_),
    .X(_1446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4536_ (.A(_1425_),
    .B_N(_1446_),
    .Y(_1447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4537_ (.B(_1446_),
    .A(_1425_),
    .X(_1448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4538_ (.A(_1441_),
    .B(_1448_),
    .Y(_1449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4539_ (.B(_1448_),
    .A(_1441_),
    .X(_1450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4540_ (.Y(_1451_),
    .A(_1428_),
    .B(_1450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4541_ (.Y(_1452_),
    .A(_1428_),
    .B(_1450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4542_ (.B(_1452_),
    .A(_1440_),
    .X(_1453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4543_ (.A(_1439_),
    .B(_1453_),
    .X(_1454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4544_ (.Y(_1455_),
    .A(_1439_),
    .B(_1453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4545_ (.A(_1455_),
    .B_N(_1438_),
    .Y(_1456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4546_ (.B(_1455_),
    .A(_1438_),
    .X(_1457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4547_ (.B1(net464),
    .VDD(VPWR),
    .Y(_1458_),
    .VSS(VGND),
    .A1(net566),
    .A2(net906));
 sg13g2_a21oi_1 _4548_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net566),
    .A2(_1457_),
    .Y(_0207_),
    .B1(_1458_));
 sg13g2_nand2_1 _4549_ (.Y(_1459_),
    .A(\mydesign.pe_weights[49] ),
    .B(\mydesign.pe_inputs[39] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4550_ (.B1(_1443_),
    .VDD(VPWR),
    .Y(_1460_),
    .VSS(VGND),
    .A1(_1442_),
    .A2(_1445_));
 sg13g2_nand2_1 _4551_ (.Y(_1461_),
    .A(\mydesign.pe_weights[50] ),
    .B(\mydesign.pe_inputs[38] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4552_ (.B(net537),
    .C(\mydesign.pe_inputs[37] ),
    .A(\mydesign.accum[68] ),
    .Y(_1462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4553_ (.A2(\mydesign.pe_inputs[37] ),
    .A1(net537),
    .B1(\mydesign.accum[68] ),
    .X(_1463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4554_ (.Y(_1464_),
    .A(_1462_),
    .B(_1463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4555_ (.B(_1464_),
    .A(_1461_),
    .X(_1465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4556_ (.Y(_1466_),
    .A(_1460_),
    .B(_1465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4557_ (.Y(_1467_),
    .A(_1460_),
    .B(_1465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4558_ (.B(_1467_),
    .A(_1459_),
    .X(_1468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4559_ (.B1(_1468_),
    .VDD(VPWR),
    .Y(_1469_),
    .VSS(VGND),
    .A1(_1447_),
    .A2(_1449_));
 sg13g2_or3_1 _4560_ (.A(_1447_),
    .B(_1449_),
    .C(_1468_),
    .X(_1470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4561_ (.A(_1469_),
    .B(_1470_),
    .X(_1471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4562_ (.B1(_1451_),
    .VDD(VPWR),
    .Y(_1472_),
    .VSS(VGND),
    .A1(_1440_),
    .A2(_1452_));
 sg13g2_nand2_1 _4563_ (.Y(_1473_),
    .A(_1471_),
    .B(_1472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4564_ (.B(_1472_),
    .A(_1471_),
    .X(_1474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4565_ (.A(_1454_),
    .B(_1456_),
    .C(_1474_),
    .X(_1475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4566_ (.B1(_1474_),
    .VDD(VPWR),
    .Y(_1476_),
    .VSS(VGND),
    .A1(_1454_),
    .A2(_1456_));
 sg13g2_a21oi_1 _4567_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1475_),
    .A2(_1476_),
    .Y(_1477_),
    .B1(net501));
 sg13g2_o21ai_1 _4568_ (.B1(net473),
    .VDD(VPWR),
    .Y(_1478_),
    .VSS(VGND),
    .A1(net574),
    .A2(net841));
 sg13g2_nor2_1 _4569_ (.A(_1477_),
    .B(_1478_),
    .Y(_0208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4570_ (.Y(_1479_),
    .A(\mydesign.pe_weights[50] ),
    .B(\mydesign.pe_inputs[39] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4571_ (.B(net537),
    .C(\mydesign.pe_inputs[38] ),
    .A(\mydesign.accum[69] ),
    .Y(_1480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4572_ (.A2(\mydesign.pe_inputs[38] ),
    .A1(net537),
    .B1(\mydesign.accum[69] ),
    .X(_1481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4573_ (.Y(_1482_),
    .A(_1480_),
    .B(_1481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4574_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1483_),
    .B(_1482_),
    .A(_1479_));
 sg13g2_xor2_1 _4575_ (.B(_1482_),
    .A(_1479_),
    .X(_1484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4576_ (.B1(_1462_),
    .VDD(VPWR),
    .Y(_1485_),
    .VSS(VGND),
    .A1(_1461_),
    .A2(_1464_));
 sg13g2_and2_1 _4577_ (.A(_1484_),
    .B(_1485_),
    .X(_1486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4578_ (.B(_1485_),
    .A(_1484_),
    .X(_1487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4579_ (.B1(_1466_),
    .VDD(VPWR),
    .Y(_1488_),
    .VSS(VGND),
    .A1(_1459_),
    .A2(_1467_));
 sg13g2_nand2_1 _4580_ (.Y(_1489_),
    .A(_1487_),
    .B(_1488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4581_ (.B(_1488_),
    .A(_1487_),
    .X(_1490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4582_ (.A(_1469_),
    .B_N(_1490_),
    .Y(_1491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4583_ (.B(_1490_),
    .A(_1469_),
    .X(_1492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4584_ (.X(_1493_),
    .A(_1473_),
    .B(_1476_),
    .C(_1492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4585_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1473_),
    .A2(_1476_),
    .Y(_1494_),
    .B1(_1492_));
 sg13g2_o21ai_1 _4586_ (.B1(net574),
    .VDD(VPWR),
    .Y(_1495_),
    .VSS(VGND),
    .A1(_1493_),
    .A2(_1494_));
 sg13g2_o21ai_1 _4587_ (.B1(net473),
    .VDD(VPWR),
    .Y(_1496_),
    .VSS(VGND),
    .A1(net574),
    .A2(net861));
 sg13g2_nor2b_1 _4588_ (.A(_1496_),
    .B_N(_1495_),
    .Y(_0209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4589_ (.B(net537),
    .C(\mydesign.pe_inputs[39] ),
    .A(\mydesign.accum[70] ),
    .Y(_1497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4590_ (.A2(\mydesign.pe_inputs[39] ),
    .A1(\mydesign.pe_weights[51] ),
    .B1(\mydesign.accum[70] ),
    .X(_1498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4591_ (.Y(_1499_),
    .A(_1497_),
    .B(_1498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4592_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1480_),
    .A2(_1483_),
    .Y(_1500_),
    .B1(_1499_));
 sg13g2_nand3_1 _4593_ (.B(_1483_),
    .C(_1499_),
    .A(_1480_),
    .Y(_1501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4594_ (.Y(_1502_),
    .B(_1501_),
    .A_N(_1500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4595_ (.Y(_1503_),
    .B(_1489_),
    .A_N(_1486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4596_ (.Y(_1504_),
    .A(_1502_),
    .B(_1503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4597_ (.A(_1491_),
    .B(_1494_),
    .C(_1504_),
    .X(_1505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4598_ (.B1(_1504_),
    .VDD(VPWR),
    .Y(_1506_),
    .VSS(VGND),
    .A1(_1491_),
    .A2(_1494_));
 sg13g2_a21oi_1 _4599_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1505_),
    .A2(_1506_),
    .Y(_1507_),
    .B1(net501));
 sg13g2_o21ai_1 _4600_ (.B1(net473),
    .VDD(VPWR),
    .Y(_1508_),
    .VSS(VGND),
    .A1(net574),
    .A2(net894));
 sg13g2_nor2_1 _4601_ (.A(_1507_),
    .B(_1508_),
    .Y(_0210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4602_ (.B1(_1506_),
    .VDD(VPWR),
    .Y(_1509_),
    .VSS(VGND),
    .A1(_1489_),
    .A2(_1502_));
 sg13g2_a21oi_1 _4603_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1486_),
    .A2(_1501_),
    .Y(_1510_),
    .B1(_1500_));
 sg13g2_xnor2_1 _4604_ (.Y(_1511_),
    .A(net843),
    .B(_1497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4605_ (.Y(_1512_),
    .A(_1510_),
    .B(_1511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4606_ (.Y(_1513_),
    .A(_1509_),
    .B(_1512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4607_ (.B1(net473),
    .VDD(VPWR),
    .Y(_1514_),
    .VSS(VGND),
    .A1(net574),
    .A2(net843));
 sg13g2_a21oi_1 _4608_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net574),
    .A2(_1513_),
    .Y(_0211_),
    .B1(_1514_));
 sg13g2_nor2_1 _4609_ (.A(net550),
    .B(\mydesign.inputs[2][16] ),
    .Y(_1515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4610_ (.A(\mydesign.inputs[2][12] ),
    .B_N(net550),
    .Y(_1516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _4611_ (.A(_0393_),
    .B(_1515_),
    .C(_1516_),
    .Y(_1517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4612_ (.A(net557),
    .B(\mydesign.inputs[2][8] ),
    .Y(_1518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4613_ (.A(\mydesign.inputs[2][4] ),
    .B_N(net557),
    .Y(_1519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4614_ (.A(_0397_),
    .B(_1518_),
    .C(_1519_),
    .Y(_1520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4615_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1521_),
    .B(_1520_),
    .A(_1517_));
 sg13g2_o21ai_1 _4616_ (.B1(net624),
    .VDD(VPWR),
    .Y(_1522_),
    .VSS(VGND),
    .A1(net485),
    .A2(_1521_));
 sg13g2_a21oi_1 _4617_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2547_),
    .A2(net492),
    .Y(_0212_),
    .B1(_1522_));
 sg13g2_mux2_1 _4618_ (.A0(\mydesign.inputs[2][17] ),
    .A1(\mydesign.inputs[2][13] ),
    .S(net550),
    .X(_1523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4619_ (.Y(_1524_),
    .A(_0392_),
    .B(_1523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4620_ (.A(net498),
    .B(\mydesign.inputs[2][5] ),
    .Y(_1525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4621_ (.B1(net460),
    .VDD(VPWR),
    .Y(_1526_),
    .VSS(VGND),
    .A1(net557),
    .A2(\mydesign.inputs[2][9] ));
 sg13g2_o21ai_1 _4622_ (.B1(_1524_),
    .VDD(VPWR),
    .Y(_1527_),
    .VSS(VGND),
    .A1(_1525_),
    .A2(_1526_));
 sg13g2_o21ai_1 _4623_ (.B1(net625),
    .VDD(VPWR),
    .Y(_1528_),
    .VSS(VGND),
    .A1(net489),
    .A2(_1527_));
 sg13g2_a21oi_1 _4624_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2546_),
    .A2(net492),
    .Y(_0213_),
    .B1(_1528_));
 sg13g2_mux2_1 _4625_ (.A0(\mydesign.inputs[2][10] ),
    .A1(\mydesign.inputs[2][6] ),
    .S(net550),
    .X(_1529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4626_ (.A0(\mydesign.inputs[2][18] ),
    .A1(\mydesign.inputs[2][14] ),
    .S(net557),
    .X(_1530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4627_ (.Y(_1531_),
    .B1(_1530_),
    .B2(_0392_),
    .A2(_1529_),
    .A1(net460),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4628_ (.B1(net625),
    .VDD(VPWR),
    .Y(_1532_),
    .VSS(VGND),
    .A1(net1090),
    .A2(net438));
 sg13g2_a21oi_1 _4629_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net438),
    .A2(_1531_),
    .Y(_0214_),
    .B1(_1532_));
 sg13g2_a21oi_1 _4630_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net557),
    .A2(_2594_),
    .Y(_1533_),
    .B1(_0397_));
 sg13g2_o21ai_1 _4631_ (.B1(_1533_),
    .VDD(VPWR),
    .Y(_1534_),
    .VSS(VGND),
    .A1(net557),
    .A2(\mydesign.inputs[2][11] ));
 sg13g2_nor2_1 _4632_ (.A(net557),
    .B(\mydesign.inputs[2][19] ),
    .Y(_1535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4633_ (.B1(_0392_),
    .VDD(VPWR),
    .Y(_1536_),
    .VSS(VGND),
    .A1(net498),
    .A2(\mydesign.inputs[2][15] ));
 sg13g2_o21ai_1 _4634_ (.B1(_1534_),
    .VDD(VPWR),
    .Y(_1537_),
    .VSS(VGND),
    .A1(_1535_),
    .A2(_1536_));
 sg13g2_o21ai_1 _4635_ (.B1(net625),
    .VDD(VPWR),
    .Y(_1538_),
    .VSS(VGND),
    .A1(net489),
    .A2(_1537_));
 sg13g2_a21oi_1 _4636_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2545_),
    .A2(net493),
    .Y(_0215_),
    .B1(_1538_));
 sg13g2_o21ai_1 _4637_ (.B1(net623),
    .VDD(VPWR),
    .Y(_1539_),
    .VSS(VGND),
    .A1(net891),
    .A2(net439));
 sg13g2_a21oi_1 _4638_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2552_),
    .A2(net439),
    .Y(_0216_),
    .B1(_1539_));
 sg13g2_o21ai_1 _4639_ (.B1(net624),
    .VDD(VPWR),
    .Y(_1540_),
    .VSS(VGND),
    .A1(\mydesign.pe_weights[29] ),
    .A2(net437));
 sg13g2_a21oi_1 _4640_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2551_),
    .A2(net437),
    .Y(_0217_),
    .B1(_1540_));
 sg13g2_o21ai_1 _4641_ (.B1(net625),
    .VDD(VPWR),
    .Y(_1541_),
    .VSS(VGND),
    .A1(\mydesign.pe_weights[30] ),
    .A2(net437));
 sg13g2_a21oi_1 _4642_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2550_),
    .A2(net437),
    .Y(_0218_),
    .B1(_1541_));
 sg13g2_o21ai_1 _4643_ (.B1(net625),
    .VDD(VPWR),
    .Y(_1542_),
    .VSS(VGND),
    .A1(net1077),
    .A2(net437));
 sg13g2_a21oi_1 _4644_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2549_),
    .A2(net437),
    .Y(_0219_),
    .B1(_1542_));
 sg13g2_and3_1 _4645_ (.X(_1543_),
    .A(net560),
    .B(\mydesign.pe_weights[44] ),
    .C(_1521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4646_ (.B1(net467),
    .VDD(VPWR),
    .Y(_1544_),
    .VSS(VGND),
    .A1(net686),
    .A2(_1543_));
 sg13g2_a21oi_1 _4647_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net686),
    .A2(_1543_),
    .Y(_0220_),
    .B1(_1544_));
 sg13g2_nand3_1 _4648_ (.B(\mydesign.pe_weights[45] ),
    .C(_1521_),
    .A(\mydesign.accum[57] ),
    .Y(_1545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4649_ (.A2(_1521_),
    .A1(\mydesign.pe_weights[45] ),
    .B1(\mydesign.accum[57] ),
    .X(_1546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4650_ (.Y(_1547_),
    .A(_1545_),
    .B(_1546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4651_ (.Y(_1548_),
    .A(\mydesign.pe_weights[44] ),
    .B(_1527_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4652_ (.A(_1547_),
    .B(_1548_),
    .Y(_1549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4653_ (.B(_1548_),
    .A(_1547_),
    .X(_1550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4654_ (.B(net815),
    .C(_1521_),
    .A(net686),
    .Y(_1551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4655_ (.B(net815),
    .C(_1521_),
    .A(net686),
    .Y(_1552_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1550_));
 sg13g2_xor2_1 _4656_ (.B(_1551_),
    .A(_1550_),
    .X(_1553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4657_ (.B1(net467),
    .VDD(VPWR),
    .Y(_1554_),
    .VSS(VGND),
    .A1(net560),
    .A2(net818));
 sg13g2_a21oi_1 _4658_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net560),
    .A2(_1553_),
    .Y(_0221_),
    .B1(_1554_));
 sg13g2_nand2b_1 _4659_ (.Y(_1555_),
    .B(\mydesign.pe_weights[44] ),
    .A_N(_1531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4660_ (.B1(\mydesign.pe_weights[46] ),
    .VDD(VPWR),
    .Y(_1556_),
    .VSS(VGND),
    .A1(_1517_),
    .A2(_1520_));
 sg13g2_nand3_1 _4661_ (.B(\mydesign.pe_weights[46] ),
    .C(_1521_),
    .A(\mydesign.accum[58] ),
    .Y(_1557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4662_ (.B(_1556_),
    .A(\mydesign.accum[58] ),
    .X(_1558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4663_ (.Y(_1559_),
    .A(\mydesign.pe_weights[45] ),
    .B(_1527_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4664_ (.A(_1558_),
    .B(_1559_),
    .Y(_1560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4665_ (.B(_1559_),
    .A(_1558_),
    .X(_1561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4666_ (.Y(_1562_),
    .B(_1561_),
    .A_N(_1545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4667_ (.Y(_1563_),
    .A(_1545_),
    .B(_1561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4668_ (.Y(_1564_),
    .B(_1563_),
    .A_N(_1555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4669_ (.Y(_1565_),
    .A(_1555_),
    .B(_1563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4670_ (.Y(_1566_),
    .A(_1549_),
    .B(_1565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4671_ (.Y(_1567_),
    .A(_1549_),
    .B(_1565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4672_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1568_),
    .B(_1567_),
    .A(_1552_));
 sg13g2_xnor2_1 _4673_ (.Y(_1569_),
    .A(_1552_),
    .B(_1567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4674_ (.B1(net467),
    .VDD(VPWR),
    .Y(_1570_),
    .VSS(VGND),
    .A1(net560),
    .A2(net959));
 sg13g2_a21oi_1 _4675_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net560),
    .A2(_1569_),
    .Y(_0222_),
    .B1(_1570_));
 sg13g2_and2_1 _4676_ (.A(_1566_),
    .B(_1568_),
    .X(_1571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4677_ (.Y(_1572_),
    .A(_1562_),
    .B(_1564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4678_ (.Y(_1573_),
    .A(\mydesign.pe_weights[44] ),
    .B(_1537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4679_ (.Y(_1574_),
    .B(\mydesign.pe_weights[45] ),
    .A_N(_1531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4680_ (.VDD(VPWR),
    .Y(_1575_),
    .A(_1574_),
    .VSS(VGND));
 sg13g2_nand2_1 _4681_ (.Y(_1576_),
    .A(\mydesign.pe_weights[46] ),
    .B(_1527_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4682_ (.B1(net535),
    .VDD(VPWR),
    .Y(_1577_),
    .VSS(VGND),
    .A1(_1517_),
    .A2(_1520_));
 sg13g2_nand3_1 _4683_ (.B(net535),
    .C(_1521_),
    .A(\mydesign.accum[59] ),
    .Y(_1578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4684_ (.A(\mydesign.accum[59] ),
    .B_N(_1577_),
    .Y(_1579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4685_ (.Y(_1580_),
    .A(\mydesign.accum[59] ),
    .B(_1577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4686_ (.Y(_1581_),
    .A(_1576_),
    .B(_1580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4687_ (.A(_1557_),
    .B_N(_1581_),
    .Y(_1582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4688_ (.Y(_1583_),
    .A(_1557_),
    .B(_1581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4689_ (.Y(_1584_),
    .A(_1574_),
    .B(_1583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4690_ (.Y(_1585_),
    .A(_1560_),
    .B(_1584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4691_ (.B(_1584_),
    .A(_1560_),
    .X(_1586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4692_ (.Y(_1587_),
    .B(_1586_),
    .A_N(_1573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4693_ (.Y(_1588_),
    .A(_1573_),
    .B(_1586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4694_ (.Y(_1589_),
    .A(_1572_),
    .B(_1588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4695_ (.Y(_1590_),
    .A(_1572_),
    .B(_1588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4696_ (.Y(_1591_),
    .A(_1571_),
    .B(_1590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4697_ (.B1(net467),
    .VDD(VPWR),
    .Y(_1592_),
    .VSS(VGND),
    .A1(net560),
    .A2(net990));
 sg13g2_a21oi_1 _4698_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net560),
    .A2(_1591_),
    .Y(_0223_),
    .B1(_1592_));
 sg13g2_o21ai_1 _4699_ (.B1(_1589_),
    .VDD(VPWR),
    .Y(_1593_),
    .VSS(VGND),
    .A1(_1571_),
    .A2(_1590_));
 sg13g2_a21oi_1 _4700_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1575_),
    .A2(_1583_),
    .Y(_1594_),
    .B1(_1582_));
 sg13g2_nand2_1 _4701_ (.Y(_1595_),
    .A(\mydesign.pe_weights[45] ),
    .B(_1537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4702_ (.B1(_1578_),
    .VDD(VPWR),
    .Y(_1596_),
    .VSS(VGND),
    .A1(_1576_),
    .A2(_1579_));
 sg13g2_nand2b_1 _4703_ (.Y(_1597_),
    .B(\mydesign.pe_weights[46] ),
    .A_N(_1531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4704_ (.B(net535),
    .C(_1527_),
    .A(\mydesign.accum[60] ),
    .Y(_1598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4705_ (.A2(_1527_),
    .A1(net535),
    .B1(\mydesign.accum[60] ),
    .X(_1599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4706_ (.Y(_1600_),
    .A(_1598_),
    .B(_1599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4707_ (.B(_1600_),
    .A(_1597_),
    .X(_1601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4708_ (.A(_1596_),
    .B(_1601_),
    .X(_1602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4709_ (.Y(_1603_),
    .A(_1596_),
    .B(_1601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4710_ (.A(_1595_),
    .B(_1603_),
    .Y(_1604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4711_ (.B(_1603_),
    .A(_1595_),
    .X(_1605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4712_ (.Y(_1606_),
    .B(_1605_),
    .A_N(_1594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4713_ (.B(_1605_),
    .A(_1594_),
    .X(_1607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4714_ (.Y(_1608_),
    .A(_1585_),
    .B(_1587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4715_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1585_),
    .A2(_1587_),
    .Y(_1609_),
    .B1(_1607_));
 sg13g2_xnor2_1 _4716_ (.Y(_1610_),
    .A(_1607_),
    .B(_1608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4717_ (.Y(_1611_),
    .A(_1593_),
    .B(_1610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4718_ (.B1(net467),
    .VDD(VPWR),
    .Y(_1612_),
    .VSS(VGND),
    .A1(net567),
    .A2(net866));
 sg13g2_a21oi_1 _4719_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net567),
    .A2(_1611_),
    .Y(_0224_),
    .B1(_1612_));
 sg13g2_a21oi_1 _4720_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1593_),
    .A2(_1610_),
    .Y(_1613_),
    .B1(_1609_));
 sg13g2_nand3b_1 _4721_ (.B(net535),
    .C(\mydesign.accum[61] ),
    .Y(_1614_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1531_));
 sg13g2_o21ai_1 _4722_ (.B1(_2548_),
    .VDD(VPWR),
    .Y(_1615_),
    .VSS(VGND),
    .A1(_2549_),
    .A2(_1531_));
 sg13g2_and2_1 _4723_ (.A(_1614_),
    .B(_1615_),
    .X(_1616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4724_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[46] ),
    .A2(_1537_),
    .Y(_1617_),
    .B1(_1616_));
 sg13g2_nand3_1 _4725_ (.B(_1537_),
    .C(_1616_),
    .A(\mydesign.pe_weights[46] ),
    .Y(_1618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4726_ (.A(_1617_),
    .B_N(_1618_),
    .Y(_1619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4727_ (.B1(_1598_),
    .VDD(VPWR),
    .Y(_1620_),
    .VSS(VGND),
    .A1(_1597_),
    .A2(_1600_));
 sg13g2_nand2_1 _4728_ (.Y(_1621_),
    .A(_1619_),
    .B(_1620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4729_ (.B(_1620_),
    .A(_1619_),
    .X(_1622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4730_ (.B1(_1622_),
    .VDD(VPWR),
    .Y(_1623_),
    .VSS(VGND),
    .A1(_1602_),
    .A2(_1604_));
 sg13g2_or3_1 _4731_ (.A(_1602_),
    .B(_1604_),
    .C(_1622_),
    .X(_1624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4732_ (.Y(_1625_),
    .A(_1623_),
    .B(_1624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4733_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1626_),
    .B(_1625_),
    .A(_1606_));
 sg13g2_xnor2_1 _4734_ (.Y(_1627_),
    .A(_1606_),
    .B(_1625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4735_ (.Y(_1628_),
    .A(_1613_),
    .B(_1627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4736_ (.B1(net469),
    .VDD(VPWR),
    .Y(_1629_),
    .VSS(VGND),
    .A1(net567),
    .A2(net840));
 sg13g2_a21oi_1 _4737_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net567),
    .A2(_1628_),
    .Y(_0225_),
    .B1(_1629_));
 sg13g2_o21ai_1 _4738_ (.B1(_1626_),
    .VDD(VPWR),
    .Y(_1630_),
    .VSS(VGND),
    .A1(_1613_),
    .A2(_1627_));
 sg13g2_a21oi_1 _4739_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net535),
    .A2(_1537_),
    .Y(_1631_),
    .B1(\mydesign.accum[62] ));
 sg13g2_nand3_1 _4740_ (.B(net535),
    .C(_1537_),
    .A(\mydesign.accum[62] ),
    .Y(_1632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4741_ (.Y(_1633_),
    .B(_1632_),
    .A_N(_1631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4742_ (.A(_1614_),
    .B(_1618_),
    .X(_1634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4743_ (.Y(_1635_),
    .A(_1633_),
    .B(_1634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4744_ (.A(_1621_),
    .B(_1635_),
    .Y(_1636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4745_ (.Y(_1637_),
    .A(_1621_),
    .B(_1635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4746_ (.A(_1623_),
    .B(_1637_),
    .Y(_1638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4747_ (.B(_1637_),
    .A(_1623_),
    .X(_1639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4748_ (.Y(_1640_),
    .A(_1630_),
    .B(_1639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4749_ (.B1(net470),
    .VDD(VPWR),
    .Y(_1641_),
    .VSS(VGND),
    .A1(net567),
    .A2(net884));
 sg13g2_a21oi_1 _4750_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net567),
    .A2(_1640_),
    .Y(_0226_),
    .B1(_1641_));
 sg13g2_a21oi_1 _4751_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1630_),
    .A2(_1639_),
    .Y(_1642_),
    .B1(_1638_));
 sg13g2_o21ai_1 _4752_ (.B1(_1632_),
    .VDD(VPWR),
    .Y(_1643_),
    .VSS(VGND),
    .A1(_1631_),
    .A2(_1634_));
 sg13g2_xor2_1 _4753_ (.B(_1643_),
    .A(net941),
    .X(_1644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4754_ (.Y(_1645_),
    .A(_1636_),
    .B(_1644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4755_ (.Y(_1646_),
    .A(_1642_),
    .B(_1645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4756_ (.B1(net470),
    .VDD(VPWR),
    .Y(_1647_),
    .VSS(VGND),
    .A1(net567),
    .A2(net941));
 sg13g2_a21oi_1 _4757_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net568),
    .A2(_1646_),
    .Y(_0227_),
    .B1(_1647_));
 sg13g2_o21ai_1 _4758_ (.B1(net637),
    .VDD(VPWR),
    .Y(_1648_),
    .VSS(VGND),
    .A1(net1022),
    .A2(net450));
 sg13g2_a21oi_1 _4759_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2547_),
    .A2(net450),
    .Y(_0228_),
    .B1(_1648_));
 sg13g2_o21ai_1 _4760_ (.B1(net637),
    .VDD(VPWR),
    .Y(_1649_),
    .VSS(VGND),
    .A1(net849),
    .A2(net447));
 sg13g2_a21oi_1 _4761_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2546_),
    .A2(net447),
    .Y(_0229_),
    .B1(_1649_));
 sg13g2_o21ai_1 _4762_ (.B1(net637),
    .VDD(VPWR),
    .Y(_1650_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[30] ),
    .A2(net493));
 sg13g2_a21oi_1 _4763_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2538_),
    .A2(net493),
    .Y(_0230_),
    .B1(_1650_));
 sg13g2_o21ai_1 _4764_ (.B1(net637),
    .VDD(VPWR),
    .Y(_1651_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[27] ),
    .A2(net447));
 sg13g2_a21oi_1 _4765_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2545_),
    .A2(net447),
    .Y(_0231_),
    .B1(_1651_));
 sg13g2_o21ai_1 _4766_ (.B1(net637),
    .VDD(VPWR),
    .Y(_1652_),
    .VSS(VGND),
    .A1(\mydesign.pe_weights[24] ),
    .A2(net451));
 sg13g2_a21oi_1 _4767_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2544_),
    .A2(net451),
    .Y(_0232_),
    .B1(_1652_));
 sg13g2_o21ai_1 _4768_ (.B1(net637),
    .VDD(VPWR),
    .Y(_1653_),
    .VSS(VGND),
    .A1(\mydesign.pe_weights[25] ),
    .A2(net451));
 sg13g2_a21oi_1 _4769_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2543_),
    .A2(net451),
    .Y(_0233_),
    .B1(_1653_));
 sg13g2_o21ai_1 _4770_ (.B1(net637),
    .VDD(VPWR),
    .Y(_1654_),
    .VSS(VGND),
    .A1(\mydesign.pe_weights[26] ),
    .A2(net452));
 sg13g2_a21oi_1 _4771_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2542_),
    .A2(net451),
    .Y(_0234_),
    .B1(_1654_));
 sg13g2_o21ai_1 _4772_ (.B1(net638),
    .VDD(VPWR),
    .Y(_1655_),
    .VSS(VGND),
    .A1(net527),
    .A2(net451));
 sg13g2_a21oi_1 _4773_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2541_),
    .A2(net451),
    .Y(_0235_),
    .B1(_1655_));
 sg13g2_nor3_1 _4774_ (.A(net502),
    .B(_2544_),
    .C(_2547_),
    .Y(_1656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4775_ (.B1(net480),
    .VDD(VPWR),
    .Y(_1657_),
    .VSS(VGND),
    .A1(net745),
    .A2(_1656_));
 sg13g2_a21oi_1 _4776_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net745),
    .A2(_1656_),
    .Y(_0236_),
    .B1(_1657_));
 sg13g2_and3_2 _4777_ (.X(_1658_),
    .A(\mydesign.accum[49] ),
    .B(\mydesign.pe_weights[41] ),
    .C(net529),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4778_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[41] ),
    .A2(net529),
    .Y(_1659_),
    .B1(\mydesign.accum[49] ));
 sg13g2_nand2_1 _4779_ (.Y(_1660_),
    .A(\mydesign.pe_weights[40] ),
    .B(\mydesign.pe_inputs[29] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4780_ (.A(_1658_),
    .B(_1659_),
    .C(_1660_),
    .Y(_1661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4781_ (.B1(_1660_),
    .VDD(VPWR),
    .Y(_1662_),
    .VSS(VGND),
    .A1(_1658_),
    .A2(_1659_));
 sg13g2_nor2b_1 _4782_ (.A(_1661_),
    .B_N(_1662_),
    .Y(_1663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4783_ (.B(\mydesign.pe_weights[40] ),
    .C(net529),
    .A(net745),
    .Y(_1664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4784_ (.B(\mydesign.pe_weights[40] ),
    .C(net529),
    .A(net745),
    .Y(_1665_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1663_));
 sg13g2_xor2_1 _4785_ (.B(_1664_),
    .A(_1663_),
    .X(_1666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4786_ (.B1(net480),
    .VDD(VPWR),
    .Y(_1667_),
    .VSS(VGND),
    .A1(net583),
    .A2(net892));
 sg13g2_a21oi_1 _4787_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net583),
    .A2(_1666_),
    .Y(_0237_),
    .B1(_1667_));
 sg13g2_nand2_1 _4788_ (.Y(_1668_),
    .A(\mydesign.pe_weights[40] ),
    .B(\mydesign.pe_inputs[30] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4789_ (.Y(_1669_),
    .A(\mydesign.pe_weights[41] ),
    .B(\mydesign.pe_inputs[29] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4790_ (.B(\mydesign.pe_weights[42] ),
    .C(net529),
    .A(\mydesign.accum[50] ),
    .Y(_1670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4791_ (.A2(net529),
    .A1(\mydesign.pe_weights[42] ),
    .B1(\mydesign.accum[50] ),
    .X(_1671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4792_ (.Y(_1672_),
    .A(_1670_),
    .B(_1671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4793_ (.A(_1669_),
    .B(_1672_),
    .Y(_1673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4794_ (.B(_1672_),
    .A(_1669_),
    .X(_1674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4795_ (.Y(_1675_),
    .A(_1658_),
    .B(_1674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4796_ (.A(_1658_),
    .B(_1674_),
    .Y(_1676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4797_ (.B(_1674_),
    .A(_1658_),
    .X(_1677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4798_ (.Y(_1678_),
    .A(_1668_),
    .B(_1677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4799_ (.Y(_1679_),
    .A(_1661_),
    .B(_1678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4800_ (.Y(_1680_),
    .A(_1661_),
    .B(_1678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4801_ (.Y(_1681_),
    .A(_1665_),
    .B(_1680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4802_ (.B1(net479),
    .VDD(VPWR),
    .Y(_1682_),
    .VSS(VGND),
    .A1(net582),
    .A2(net900));
 sg13g2_a21oi_1 _4803_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net582),
    .A2(_1681_),
    .Y(_0238_),
    .B1(_1682_));
 sg13g2_o21ai_1 _4804_ (.B1(_1679_),
    .VDD(VPWR),
    .Y(_1683_),
    .VSS(VGND),
    .A1(_1665_),
    .A2(_1680_));
 sg13g2_o21ai_1 _4805_ (.B1(_1675_),
    .VDD(VPWR),
    .Y(_1684_),
    .VSS(VGND),
    .A1(_1668_),
    .A2(_1676_));
 sg13g2_nand2_1 _4806_ (.Y(_1685_),
    .A(\mydesign.pe_weights[40] ),
    .B(\mydesign.pe_inputs[31] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4807_ (.Y(_1686_),
    .A(\mydesign.pe_weights[41] ),
    .B(\mydesign.pe_inputs[30] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4808_ (.Y(_1687_),
    .A(\mydesign.pe_weights[42] ),
    .B(\mydesign.pe_inputs[29] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4809_ (.B(net533),
    .C(net529),
    .A(\mydesign.accum[51] ),
    .Y(_1688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4810_ (.A2(\mydesign.pe_inputs[28] ),
    .A1(net533),
    .B1(\mydesign.accum[51] ),
    .X(_1689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4811_ (.Y(_1690_),
    .A(_1688_),
    .B(_1689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4812_ (.B(_1690_),
    .A(_1687_),
    .X(_1691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4813_ (.A(_1670_),
    .B_N(_1691_),
    .Y(_1692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4814_ (.B(_1691_),
    .A(_1670_),
    .X(_1693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4815_ (.A(_1686_),
    .B(_1693_),
    .Y(_1694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4816_ (.B(_1693_),
    .A(_1686_),
    .X(_1695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4817_ (.Y(_1696_),
    .A(_1673_),
    .B(_1695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4818_ (.Y(_1697_),
    .A(_1673_),
    .B(_1695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4819_ (.B(_1697_),
    .A(_1685_),
    .X(_1698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4820_ (.A(_1684_),
    .B(_1698_),
    .X(_1699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4821_ (.Y(_1700_),
    .A(_1684_),
    .B(_1698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4822_ (.A(_1700_),
    .B_N(_1683_),
    .Y(_1701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4823_ (.B(_1700_),
    .A(_1683_),
    .X(_1702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4824_ (.B1(net479),
    .VDD(VPWR),
    .Y(_1703_),
    .VSS(VGND),
    .A1(net582),
    .A2(net969));
 sg13g2_a21oi_1 _4825_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net582),
    .A2(_1702_),
    .Y(_0239_),
    .B1(_1703_));
 sg13g2_nand2_1 _4826_ (.Y(_1704_),
    .A(\mydesign.pe_weights[41] ),
    .B(\mydesign.pe_inputs[31] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4827_ (.B1(_1688_),
    .VDD(VPWR),
    .Y(_1705_),
    .VSS(VGND),
    .A1(_1687_),
    .A2(_1690_));
 sg13g2_nand2_1 _4828_ (.Y(_1706_),
    .A(\mydesign.pe_weights[42] ),
    .B(\mydesign.pe_inputs[30] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4829_ (.B(net533),
    .C(\mydesign.pe_inputs[29] ),
    .A(\mydesign.accum[52] ),
    .Y(_1707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4830_ (.A2(\mydesign.pe_inputs[29] ),
    .A1(net533),
    .B1(\mydesign.accum[52] ),
    .X(_1708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4831_ (.Y(_1709_),
    .A(_1707_),
    .B(_1708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4832_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1710_),
    .B(_1709_),
    .A(_1706_));
 sg13g2_xor2_1 _4833_ (.B(_1709_),
    .A(_1706_),
    .X(_1711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4834_ (.Y(_1712_),
    .A(_1705_),
    .B(_1711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4835_ (.Y(_1713_),
    .A(_1705_),
    .B(_1711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4836_ (.B(_1713_),
    .A(_1704_),
    .X(_1714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4837_ (.B1(_1714_),
    .VDD(VPWR),
    .Y(_1715_),
    .VSS(VGND),
    .A1(_1692_),
    .A2(_1694_));
 sg13g2_or3_1 _4838_ (.A(_1692_),
    .B(_1694_),
    .C(_1714_),
    .X(_1716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4839_ (.A(_1715_),
    .B(_1716_),
    .X(_1717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4840_ (.B1(_1696_),
    .VDD(VPWR),
    .Y(_1718_),
    .VSS(VGND),
    .A1(_1685_),
    .A2(_1697_));
 sg13g2_nand2_1 _4841_ (.Y(_1719_),
    .A(_1717_),
    .B(_1718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4842_ (.B(_1718_),
    .A(_1717_),
    .X(_1720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4843_ (.A(_1699_),
    .B(_1701_),
    .C(_1720_),
    .X(_1721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4844_ (.B1(_1720_),
    .VDD(VPWR),
    .Y(_1722_),
    .VSS(VGND),
    .A1(_1699_),
    .A2(_1701_));
 sg13g2_a21oi_1 _4845_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1721_),
    .A2(_1722_),
    .Y(_1723_),
    .B1(net502));
 sg13g2_o21ai_1 _4846_ (.B1(net479),
    .VDD(VPWR),
    .Y(_1724_),
    .VSS(VGND),
    .A1(net582),
    .A2(net926));
 sg13g2_nor2_1 _4847_ (.A(_1723_),
    .B(_1724_),
    .Y(_0240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4848_ (.B1(_1712_),
    .VDD(VPWR),
    .Y(_1725_),
    .VSS(VGND),
    .A1(_1704_),
    .A2(_1713_));
 sg13g2_nand2_1 _4849_ (.Y(_1726_),
    .A(\mydesign.pe_weights[42] ),
    .B(\mydesign.pe_inputs[31] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4850_ (.B(net533),
    .C(\mydesign.pe_inputs[30] ),
    .A(\mydesign.accum[53] ),
    .Y(_1727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4851_ (.A2(\mydesign.pe_inputs[30] ),
    .A1(net533),
    .B1(\mydesign.accum[53] ),
    .X(_1728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4852_ (.Y(_1729_),
    .A(_1727_),
    .B(_1728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4853_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1730_),
    .B(_1729_),
    .A(_1726_));
 sg13g2_xnor2_1 _4854_ (.Y(_1731_),
    .A(_1726_),
    .B(_1729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4855_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1707_),
    .A2(_1710_),
    .Y(_1732_),
    .B1(_1731_));
 sg13g2_nand3_1 _4856_ (.B(_1710_),
    .C(_1731_),
    .A(_1707_),
    .Y(_1733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4857_ (.A(_1732_),
    .B_N(_1733_),
    .Y(_1734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4858_ (.Y(_1735_),
    .A(_1725_),
    .B(_1734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4859_ (.Y(_1736_),
    .A(_1725_),
    .B(_1734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4860_ (.A(_1715_),
    .B(_1736_),
    .Y(_1737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4861_ (.Y(_1738_),
    .A(_1715_),
    .B(_1736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4862_ (.X(_1739_),
    .A(_1719_),
    .B(_1722_),
    .C(_1738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4863_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1719_),
    .A2(_1722_),
    .Y(_1740_),
    .B1(_1738_));
 sg13g2_o21ai_1 _4864_ (.B1(net582),
    .VDD(VPWR),
    .Y(_1741_),
    .VSS(VGND),
    .A1(_1739_),
    .A2(_1740_));
 sg13g2_o21ai_1 _4865_ (.B1(net479),
    .VDD(VPWR),
    .Y(_1742_),
    .VSS(VGND),
    .A1(net582),
    .A2(net918));
 sg13g2_nor2b_1 _4866_ (.A(_1742_),
    .B_N(_1741_),
    .Y(_0241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4867_ (.B(net533),
    .C(\mydesign.pe_inputs[31] ),
    .A(\mydesign.accum[54] ),
    .Y(_1743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4868_ (.A2(\mydesign.pe_inputs[31] ),
    .A1(\mydesign.pe_weights[43] ),
    .B1(\mydesign.accum[54] ),
    .X(_1744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4869_ (.Y(_1745_),
    .A(_1743_),
    .B(_1744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4870_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1727_),
    .A2(_1730_),
    .Y(_1746_),
    .B1(_1745_));
 sg13g2_nand3_1 _4871_ (.B(_1730_),
    .C(_1745_),
    .A(_1727_),
    .Y(_1747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4872_ (.Y(_1748_),
    .B(_1747_),
    .A_N(_1746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4873_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1725_),
    .A2(_1733_),
    .Y(_1749_),
    .B1(_1732_));
 sg13g2_xor2_1 _4874_ (.B(_1749_),
    .A(_1748_),
    .X(_1750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4875_ (.A(_1737_),
    .B(_1740_),
    .C(_1750_),
    .X(_1751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4876_ (.B1(_1750_),
    .VDD(VPWR),
    .Y(_1752_),
    .VSS(VGND),
    .A1(_1737_),
    .A2(_1740_));
 sg13g2_a21oi_1 _4877_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1751_),
    .A2(_1752_),
    .Y(_1753_),
    .B1(net502));
 sg13g2_o21ai_1 _4878_ (.B1(net482),
    .VDD(VPWR),
    .Y(_1754_),
    .VSS(VGND),
    .A1(net582),
    .A2(net827));
 sg13g2_nor2_1 _4879_ (.A(_1753_),
    .B(_1754_),
    .Y(_0242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4880_ (.B1(_1752_),
    .VDD(VPWR),
    .Y(_1755_),
    .VSS(VGND),
    .A1(_1735_),
    .A2(_1748_));
 sg13g2_a21oi_1 _4881_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1732_),
    .A2(_1747_),
    .Y(_1756_),
    .B1(_1746_));
 sg13g2_xnor2_1 _4882_ (.Y(_1757_),
    .A(net912),
    .B(_1743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4883_ (.Y(_1758_),
    .A(_1756_),
    .B(_1757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4884_ (.Y(_1759_),
    .A(_1755_),
    .B(_1758_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4885_ (.B1(net479),
    .VDD(VPWR),
    .Y(_1760_),
    .VSS(VGND),
    .A1(net590),
    .A2(net912));
 sg13g2_a21oi_1 _4886_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net583),
    .A2(_1759_),
    .Y(_0243_),
    .B1(_1760_));
 sg13g2_or3_1 _4887_ (.A(_2606_),
    .B(_2607_),
    .C(_2618_),
    .X(_1761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4888_ (.A(net623),
    .B(_1761_),
    .X(_1762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4889_ (.Y(_1763_),
    .A(net654),
    .B(_1762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4890_ (.B1(_1763_),
    .VDD(VPWR),
    .Y(_0244_),
    .VSS(VGND),
    .A1(net603),
    .A2(_1761_));
 sg13g2_nand2_1 _4891_ (.Y(_1764_),
    .A(net697),
    .B(_1762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4892_ (.B1(_1764_),
    .VDD(VPWR),
    .Y(_0245_),
    .VSS(VGND),
    .A1(net601),
    .A2(_1761_));
 sg13g2_nand2_1 _4893_ (.Y(_1765_),
    .A(net671),
    .B(_1762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4894_ (.B1(_1765_),
    .VDD(VPWR),
    .Y(_0246_),
    .VSS(VGND),
    .A1(net599),
    .A2(_1761_));
 sg13g2_nand2_1 _4895_ (.Y(_1766_),
    .A(net648),
    .B(_1762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4896_ (.B1(_1766_),
    .VDD(VPWR),
    .Y(_0247_),
    .VSS(VGND),
    .A1(net597),
    .A2(_1761_));
 sg13g2_nor3_2 _4897_ (.A(_2591_),
    .B(_2648_),
    .C(_2657_),
    .Y(_1767_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _4898_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2605_),
    .Y(_1768_),
    .A2(_2688_),
    .A1(_2664_));
 sg13g2_nand2_2 _4899_ (.Y(_1769_),
    .A(net1),
    .B(_1768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4900_ (.B1(net612),
    .VDD(VPWR),
    .Y(_1770_),
    .VSS(VGND),
    .A1(net844),
    .A2(_1767_));
 sg13g2_a21oi_1 _4901_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1767_),
    .A2(_1769_),
    .Y(_0248_),
    .B1(net845));
 sg13g2_nand2_2 _4902_ (.Y(_1771_),
    .A(net2),
    .B(_1768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4903_ (.B1(net612),
    .VDD(VPWR),
    .Y(_1772_),
    .VSS(VGND),
    .A1(net858),
    .A2(_1767_));
 sg13g2_a21oi_1 _4904_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1767_),
    .A2(_1771_),
    .Y(_0249_),
    .B1(net859));
 sg13g2_nand2_2 _4905_ (.Y(_1773_),
    .A(net3),
    .B(_1768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4906_ (.B1(net613),
    .VDD(VPWR),
    .Y(_1774_),
    .VSS(VGND),
    .A1(net853),
    .A2(_1767_));
 sg13g2_a21oi_1 _4907_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1767_),
    .A2(_1773_),
    .Y(_0250_),
    .B1(net854));
 sg13g2_nand2_1 _4908_ (.Y(_1775_),
    .A(net4),
    .B(_1768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4909_ (.B1(net612),
    .VDD(VPWR),
    .Y(_1776_),
    .VSS(VGND),
    .A1(net820),
    .A2(_1767_));
 sg13g2_a21oi_1 _4910_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1767_),
    .A2(_1775_),
    .Y(_0251_),
    .B1(net821));
 sg13g2_o21ai_1 _4911_ (.B1(net634),
    .VDD(VPWR),
    .Y(_1777_),
    .VSS(VGND),
    .A1(net526),
    .A2(net442));
 sg13g2_a21oi_1 _4912_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2540_),
    .A2(net442),
    .Y(_0252_),
    .B1(_1777_));
 sg13g2_o21ai_1 _4913_ (.B1(net634),
    .VDD(VPWR),
    .Y(_1778_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[21] ),
    .A2(net442));
 sg13g2_a21oi_1 _4914_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2539_),
    .A2(net442),
    .Y(_0253_),
    .B1(_1778_));
 sg13g2_o21ai_1 _4915_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1779_),
    .VSS(VGND),
    .A1(net1037),
    .A2(net442));
 sg13g2_a21oi_1 _4916_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2538_),
    .A2(net442),
    .Y(_0254_),
    .B1(_1779_));
 sg13g2_o21ai_1 _4917_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1780_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[23] ),
    .A2(net440));
 sg13g2_a21oi_1 _4918_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2537_),
    .A2(net440),
    .Y(_0255_),
    .B1(_1780_));
 sg13g2_o21ai_1 _4919_ (.B1(net635),
    .VDD(VPWR),
    .Y(_1781_),
    .VSS(VGND),
    .A1(net1043),
    .A2(net444));
 sg13g2_a21oi_1 _4920_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2536_),
    .A2(net445),
    .Y(_0256_),
    .B1(_1781_));
 sg13g2_o21ai_1 _4921_ (.B1(net635),
    .VDD(VPWR),
    .Y(_1782_),
    .VSS(VGND),
    .A1(\mydesign.pe_weights[21] ),
    .A2(net445));
 sg13g2_a21oi_1 _4922_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2535_),
    .A2(net445),
    .Y(_0257_),
    .B1(_1782_));
 sg13g2_o21ai_1 _4923_ (.B1(net638),
    .VDD(VPWR),
    .Y(_1783_),
    .VSS(VGND),
    .A1(net525),
    .A2(net449));
 sg13g2_a21oi_1 _4924_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2534_),
    .A2(net449),
    .Y(_0258_),
    .B1(_1783_));
 sg13g2_o21ai_1 _4925_ (.B1(net638),
    .VDD(VPWR),
    .Y(_1784_),
    .VSS(VGND),
    .A1(net1025),
    .A2(net449));
 sg13g2_a21oi_1 _4926_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2533_),
    .A2(net449),
    .Y(_0259_),
    .B1(_1784_));
 sg13g2_nor3_1 _4927_ (.A(net501),
    .B(_2536_),
    .C(_2540_),
    .Y(_1785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4928_ (.B1(net477),
    .VDD(VPWR),
    .Y(_1786_),
    .VSS(VGND),
    .A1(net664),
    .A2(_1785_));
 sg13g2_a21oi_1 _4929_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net664),
    .A2(_1785_),
    .Y(_0260_),
    .B1(_1786_));
 sg13g2_and3_2 _4930_ (.X(_1787_),
    .A(\mydesign.accum[41] ),
    .B(\mydesign.pe_weights[37] ),
    .C(net528),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4931_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[37] ),
    .A2(net528),
    .Y(_1788_),
    .B1(\mydesign.accum[41] ));
 sg13g2_nand2_1 _4932_ (.Y(_1789_),
    .A(\mydesign.pe_weights[36] ),
    .B(\mydesign.pe_inputs[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4933_ (.A(_1787_),
    .B(_1788_),
    .C(_1789_),
    .Y(_1790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4934_ (.B1(_1789_),
    .VDD(VPWR),
    .Y(_1791_),
    .VSS(VGND),
    .A1(_1787_),
    .A2(_1788_));
 sg13g2_nor2b_1 _4935_ (.A(_1790_),
    .B_N(_1791_),
    .Y(_1792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4936_ (.B(net943),
    .C(net528),
    .A(net664),
    .Y(_1793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4937_ (.B(\mydesign.pe_weights[36] ),
    .C(net528),
    .A(net664),
    .Y(_1794_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1792_));
 sg13g2_xor2_1 _4938_ (.B(_1793_),
    .A(_1792_),
    .X(_1795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4939_ (.B1(net477),
    .VDD(VPWR),
    .Y(_1796_),
    .VSS(VGND),
    .A1(net585),
    .A2(net949));
 sg13g2_a21oi_1 _4940_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net585),
    .A2(_1795_),
    .Y(_0261_),
    .B1(_1796_));
 sg13g2_nand2_1 _4941_ (.Y(_1797_),
    .A(\mydesign.pe_weights[36] ),
    .B(\mydesign.pe_inputs[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4942_ (.Y(_1798_),
    .A(\mydesign.pe_weights[37] ),
    .B(\mydesign.pe_inputs[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4943_ (.B(\mydesign.pe_weights[38] ),
    .C(net528),
    .A(\mydesign.accum[42] ),
    .Y(_1799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4944_ (.A2(net528),
    .A1(\mydesign.pe_weights[38] ),
    .B1(\mydesign.accum[42] ),
    .X(_1800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4945_ (.Y(_1801_),
    .A(_1799_),
    .B(_1800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4946_ (.A(_1798_),
    .B(_1801_),
    .Y(_1802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4947_ (.B(_1801_),
    .A(_1798_),
    .X(_1803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4948_ (.Y(_1804_),
    .A(_1787_),
    .B(_1803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4949_ (.A(_1787_),
    .B(_1803_),
    .Y(_1805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4950_ (.B(_1803_),
    .A(_1787_),
    .X(_1806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4951_ (.Y(_1807_),
    .A(_1797_),
    .B(_1806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4952_ (.Y(_1808_),
    .A(_1790_),
    .B(_1807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4953_ (.Y(_1809_),
    .A(_1790_),
    .B(_1807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4954_ (.Y(_1810_),
    .A(_1794_),
    .B(_1809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4955_ (.B1(net478),
    .VDD(VPWR),
    .Y(_1811_),
    .VSS(VGND),
    .A1(net589),
    .A2(net921));
 sg13g2_a21oi_1 _4956_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net589),
    .A2(_1810_),
    .Y(_0262_),
    .B1(_1811_));
 sg13g2_o21ai_1 _4957_ (.B1(_1808_),
    .VDD(VPWR),
    .Y(_1812_),
    .VSS(VGND),
    .A1(_1794_),
    .A2(_1809_));
 sg13g2_o21ai_1 _4958_ (.B1(_1804_),
    .VDD(VPWR),
    .Y(_1813_),
    .VSS(VGND),
    .A1(_1797_),
    .A2(_1805_));
 sg13g2_nand2_1 _4959_ (.Y(_1814_),
    .A(\mydesign.pe_weights[36] ),
    .B(\mydesign.pe_inputs[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4960_ (.Y(_1815_),
    .A(\mydesign.pe_weights[37] ),
    .B(\mydesign.pe_inputs[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4961_ (.Y(_1816_),
    .A(\mydesign.pe_weights[38] ),
    .B(\mydesign.pe_inputs[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4962_ (.B(net531),
    .C(net528),
    .A(\mydesign.accum[43] ),
    .Y(_1817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4963_ (.A2(\mydesign.pe_inputs[24] ),
    .A1(net531),
    .B1(\mydesign.accum[43] ),
    .X(_1818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4964_ (.Y(_1819_),
    .A(_1817_),
    .B(_1818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4965_ (.B(_1819_),
    .A(_1816_),
    .X(_1820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4966_ (.A(_1799_),
    .B_N(_1820_),
    .Y(_1821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4967_ (.B(_1820_),
    .A(_1799_),
    .X(_1822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4968_ (.A(_1815_),
    .B(_1822_),
    .Y(_1823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4969_ (.B(_1822_),
    .A(_1815_),
    .X(_1824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4970_ (.Y(_1825_),
    .A(_1802_),
    .B(_1824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4971_ (.Y(_1826_),
    .A(_1802_),
    .B(_1824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4972_ (.B(_1826_),
    .A(_1814_),
    .X(_1827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4973_ (.A(_1813_),
    .B(_1827_),
    .X(_1828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4974_ (.Y(_1829_),
    .A(_1813_),
    .B(_1827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4975_ (.A(_1829_),
    .B_N(_1812_),
    .Y(_1830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4976_ (.B(_1829_),
    .A(_1812_),
    .X(_1831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4977_ (.B1(net474),
    .VDD(VPWR),
    .Y(_1832_),
    .VSS(VGND),
    .A1(net585),
    .A2(net902));
 sg13g2_a21oi_1 _4978_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net585),
    .A2(_1831_),
    .Y(_0263_),
    .B1(_1832_));
 sg13g2_nand2_1 _4979_ (.Y(_1833_),
    .A(\mydesign.pe_weights[37] ),
    .B(\mydesign.pe_inputs[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4980_ (.B1(_1817_),
    .VDD(VPWR),
    .Y(_1834_),
    .VSS(VGND),
    .A1(_1816_),
    .A2(_1819_));
 sg13g2_nand2_1 _4981_ (.Y(_1835_),
    .A(\mydesign.pe_weights[38] ),
    .B(\mydesign.pe_inputs[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4982_ (.B(net531),
    .C(\mydesign.pe_inputs[25] ),
    .A(\mydesign.accum[44] ),
    .Y(_1836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4983_ (.A2(\mydesign.pe_inputs[25] ),
    .A1(net531),
    .B1(\mydesign.accum[44] ),
    .X(_1837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4984_ (.Y(_1838_),
    .A(_1836_),
    .B(_1837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4985_ (.B(_1838_),
    .A(_1835_),
    .X(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4986_ (.A(_1834_),
    .B(_1839_),
    .X(_1840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4987_ (.Y(_1841_),
    .A(_1834_),
    .B(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4988_ (.A(_1833_),
    .B(_1841_),
    .Y(_1842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4989_ (.B(_1841_),
    .A(_1833_),
    .X(_1843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4990_ (.B1(_1843_),
    .VDD(VPWR),
    .Y(_1844_),
    .VSS(VGND),
    .A1(_1821_),
    .A2(_1823_));
 sg13g2_or3_1 _4991_ (.A(_1821_),
    .B(_1823_),
    .C(_1843_),
    .X(_1845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4992_ (.A(_1844_),
    .B(_1845_),
    .X(_1846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4993_ (.B1(_1825_),
    .VDD(VPWR),
    .Y(_1847_),
    .VSS(VGND),
    .A1(_1814_),
    .A2(_1826_));
 sg13g2_nand2_1 _4994_ (.Y(_1848_),
    .A(_1846_),
    .B(_1847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4995_ (.B(_1847_),
    .A(_1846_),
    .X(_1849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4996_ (.A(_1828_),
    .B(_1830_),
    .C(_1849_),
    .X(_1850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4997_ (.B1(_1849_),
    .VDD(VPWR),
    .Y(_1851_),
    .VSS(VGND),
    .A1(_1828_),
    .A2(_1830_));
 sg13g2_a21oi_1 _4998_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1850_),
    .A2(_1851_),
    .Y(_1852_),
    .B1(net501));
 sg13g2_o21ai_1 _4999_ (.B1(net477),
    .VDD(VPWR),
    .Y(_1853_),
    .VSS(VGND),
    .A1(net585),
    .A2(net1018));
 sg13g2_nor2_1 _5000_ (.A(_1852_),
    .B(_1853_),
    .Y(_0264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5001_ (.Y(_1854_),
    .A(\mydesign.pe_weights[38] ),
    .B(\mydesign.pe_inputs[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5002_ (.B(net531),
    .C(\mydesign.pe_inputs[26] ),
    .A(\mydesign.accum[45] ),
    .Y(_1855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5003_ (.A2(\mydesign.pe_inputs[26] ),
    .A1(net531),
    .B1(\mydesign.accum[45] ),
    .X(_1856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5004_ (.Y(_1857_),
    .A(_1855_),
    .B(_1856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5005_ (.B(_1857_),
    .A(_1854_),
    .X(_1858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5006_ (.B1(_1836_),
    .VDD(VPWR),
    .Y(_1859_),
    .VSS(VGND),
    .A1(_1835_),
    .A2(_1838_));
 sg13g2_nand2_1 _5007_ (.Y(_1860_),
    .A(_1858_),
    .B(_1859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5008_ (.B(_1859_),
    .A(_1858_),
    .X(_1861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5009_ (.B1(_1861_),
    .VDD(VPWR),
    .Y(_1862_),
    .VSS(VGND),
    .A1(_1840_),
    .A2(_1842_));
 sg13g2_or3_1 _5010_ (.A(_1840_),
    .B(_1842_),
    .C(_1861_),
    .X(_1863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5011_ (.A(_1862_),
    .B(_1863_),
    .X(_1864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5012_ (.A(_1844_),
    .B_N(_1864_),
    .Y(_1865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5013_ (.B(_1864_),
    .A(_1844_),
    .X(_1866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5014_ (.X(_1867_),
    .A(_1848_),
    .B(_1851_),
    .C(_1866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5015_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1848_),
    .A2(_1851_),
    .Y(_1868_),
    .B1(_1866_));
 sg13g2_o21ai_1 _5016_ (.B1(net591),
    .VDD(VPWR),
    .Y(_1869_),
    .VSS(VGND),
    .A1(_1867_),
    .A2(_1868_));
 sg13g2_o21ai_1 _5017_ (.B1(_1869_),
    .VDD(VPWR),
    .Y(_1870_),
    .VSS(VGND),
    .A1(net591),
    .A2(net1019));
 sg13g2_nor2_1 _5018_ (.A(net463),
    .B(_1870_),
    .Y(_0265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5019_ (.Y(_1871_),
    .A(_1860_),
    .B(_1862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5020_ (.B(net531),
    .C(\mydesign.pe_inputs[27] ),
    .A(\mydesign.accum[46] ),
    .Y(_1872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5021_ (.A2(\mydesign.pe_inputs[27] ),
    .A1(\mydesign.pe_weights[39] ),
    .B1(\mydesign.accum[46] ),
    .X(_1873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5022_ (.Y(_1874_),
    .A(_1872_),
    .B(_1873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5023_ (.B1(_1855_),
    .VDD(VPWR),
    .Y(_1875_),
    .VSS(VGND),
    .A1(_1854_),
    .A2(_1857_));
 sg13g2_nor2b_1 _5024_ (.A(_1875_),
    .B_N(_1874_),
    .Y(_1876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5025_ (.Y(_1877_),
    .B(_1875_),
    .A_N(_1874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5026_ (.Y(_1878_),
    .B(_1877_),
    .A_N(_1876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5027_ (.Y(_1879_),
    .A(_1871_),
    .B(_1878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5028_ (.A(_1865_),
    .B(_1868_),
    .C(_1879_),
    .X(_1880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5029_ (.B1(_1879_),
    .VDD(VPWR),
    .Y(_1881_),
    .VSS(VGND),
    .A1(_1865_),
    .A2(_1868_));
 sg13g2_a21oi_1 _5030_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1880_),
    .A2(_1881_),
    .Y(_1882_),
    .B1(net502));
 sg13g2_o21ai_1 _5031_ (.B1(net480),
    .VDD(VPWR),
    .Y(_1883_),
    .VSS(VGND),
    .A1(net591),
    .A2(net963));
 sg13g2_nor2_1 _5032_ (.A(_1882_),
    .B(_1883_),
    .Y(_0266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5033_ (.B1(_1881_),
    .VDD(VPWR),
    .Y(_1884_),
    .VSS(VGND),
    .A1(_1862_),
    .A2(_1878_));
 sg13g2_a21oi_1 _5034_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1860_),
    .A2(_1877_),
    .Y(_1885_),
    .B1(_1876_));
 sg13g2_xor2_1 _5035_ (.B(_1872_),
    .A(net980),
    .X(_1886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5036_ (.Y(_1887_),
    .A(_1885_),
    .B(_1886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5037_ (.Y(_1888_),
    .A(_1884_),
    .B(_1887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5038_ (.B1(net480),
    .VDD(VPWR),
    .Y(_1889_),
    .VSS(VGND),
    .A1(net583),
    .A2(net980));
 sg13g2_a21oi_1 _5039_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net583),
    .A2(_1888_),
    .Y(_0267_),
    .B1(_1889_));
 sg13g2_o21ai_1 _5040_ (.B1(net634),
    .VDD(VPWR),
    .Y(_1890_),
    .VSS(VGND),
    .A1(net903),
    .A2(net443));
 sg13g2_a21oi_1 _5041_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2532_),
    .A2(net443),
    .Y(_0268_),
    .B1(_1890_));
 sg13g2_o21ai_1 _5042_ (.B1(net634),
    .VDD(VPWR),
    .Y(_1891_),
    .VSS(VGND),
    .A1(\mydesign.pe_weights[17] ),
    .A2(net443));
 sg13g2_a21oi_1 _5043_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2531_),
    .A2(net443),
    .Y(_0269_),
    .B1(_1891_));
 sg13g2_o21ai_1 _5044_ (.B1(net634),
    .VDD(VPWR),
    .Y(_1892_),
    .VSS(VGND),
    .A1(net1017),
    .A2(net443));
 sg13g2_a21oi_1 _5045_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2530_),
    .A2(net442),
    .Y(_0270_),
    .B1(_1892_));
 sg13g2_o21ai_1 _5046_ (.B1(net634),
    .VDD(VPWR),
    .Y(_1893_),
    .VSS(VGND),
    .A1(\mydesign.pe_weights[19] ),
    .A2(net442));
 sg13g2_a21oi_1 _5047_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2529_),
    .A2(net443),
    .Y(_0271_),
    .B1(_1893_));
 sg13g2_and3_1 _5048_ (.X(_1894_),
    .A(net584),
    .B(\mydesign.pe_weights[32] ),
    .C(net526),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5049_ (.B1(net475),
    .VDD(VPWR),
    .Y(_1895_),
    .VSS(VGND),
    .A1(net734),
    .A2(_1894_));
 sg13g2_a21oi_1 _5050_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net734),
    .A2(_1894_),
    .Y(_0272_),
    .B1(_1895_));
 sg13g2_and3_2 _5051_ (.X(_1896_),
    .A(\mydesign.accum[33] ),
    .B(\mydesign.pe_weights[33] ),
    .C(net526),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5052_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[33] ),
    .A2(net526),
    .Y(_1897_),
    .B1(\mydesign.accum[33] ));
 sg13g2_nand2_1 _5053_ (.Y(_1898_),
    .A(\mydesign.pe_weights[32] ),
    .B(\mydesign.pe_inputs[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5054_ (.A(_1896_),
    .B(_1897_),
    .C(_1898_),
    .Y(_1899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5055_ (.B1(_1898_),
    .VDD(VPWR),
    .Y(_1900_),
    .VSS(VGND),
    .A1(_1896_),
    .A2(_1897_));
 sg13g2_nor2b_1 _5056_ (.A(_1899_),
    .B_N(_1900_),
    .Y(_1901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5057_ (.B(\mydesign.pe_weights[32] ),
    .C(net526),
    .A(net734),
    .Y(_1902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5058_ (.B(\mydesign.pe_weights[32] ),
    .C(net1107),
    .A(net734),
    .Y(_1903_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1901_));
 sg13g2_xor2_1 _5059_ (.B(_1902_),
    .A(_1901_),
    .X(_1904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5060_ (.B1(net475),
    .VDD(VPWR),
    .Y(_1905_),
    .VSS(VGND),
    .A1(net584),
    .A2(net919));
 sg13g2_a21oi_1 _5061_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net584),
    .A2(_1904_),
    .Y(_0273_),
    .B1(_1905_));
 sg13g2_nand2_1 _5062_ (.Y(_1906_),
    .A(\mydesign.pe_weights[32] ),
    .B(\mydesign.pe_inputs[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5063_ (.Y(_1907_),
    .A(\mydesign.pe_weights[33] ),
    .B(\mydesign.pe_inputs[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5064_ (.B(net530),
    .C(net526),
    .A(\mydesign.accum[34] ),
    .Y(_1908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5065_ (.A2(net526),
    .A1(net530),
    .B1(\mydesign.accum[34] ),
    .X(_1909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5066_ (.Y(_1910_),
    .A(_1908_),
    .B(_1909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5067_ (.A(_1907_),
    .B(_1910_),
    .Y(_1911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5068_ (.B(_1910_),
    .A(_1907_),
    .X(_1912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5069_ (.Y(_1913_),
    .A(_1896_),
    .B(_1912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5070_ (.A(_1896_),
    .B(_1912_),
    .Y(_1914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5071_ (.B(_1912_),
    .A(_1896_),
    .X(_1915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5072_ (.Y(_1916_),
    .A(_1906_),
    .B(_1915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5073_ (.Y(_1917_),
    .A(_1899_),
    .B(_1916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5074_ (.Y(_1918_),
    .A(_1899_),
    .B(_1916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5075_ (.Y(_1919_),
    .A(_1903_),
    .B(_1918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5076_ (.B1(net475),
    .VDD(VPWR),
    .Y(_1920_),
    .VSS(VGND),
    .A1(net584),
    .A2(net913));
 sg13g2_a21oi_1 _5077_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net584),
    .A2(_1919_),
    .Y(_0274_),
    .B1(_1920_));
 sg13g2_o21ai_1 _5078_ (.B1(_1917_),
    .VDD(VPWR),
    .Y(_1921_),
    .VSS(VGND),
    .A1(_1903_),
    .A2(_1918_));
 sg13g2_o21ai_1 _5079_ (.B1(_1913_),
    .VDD(VPWR),
    .Y(_1922_),
    .VSS(VGND),
    .A1(_1906_),
    .A2(_1914_));
 sg13g2_nand2_1 _5080_ (.Y(_1923_),
    .A(\mydesign.pe_weights[32] ),
    .B(\mydesign.pe_inputs[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5081_ (.Y(_1924_),
    .A(\mydesign.pe_weights[33] ),
    .B(\mydesign.pe_inputs[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5082_ (.Y(_1925_),
    .A(\mydesign.pe_weights[35] ),
    .B(net526),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5083_ (.B(\mydesign.pe_weights[34] ),
    .C(\mydesign.pe_inputs[21] ),
    .A(\mydesign.accum[35] ),
    .Y(_1926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5084_ (.A2(\mydesign.pe_inputs[21] ),
    .A1(\mydesign.pe_weights[34] ),
    .B1(\mydesign.accum[35] ),
    .X(_1927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5085_ (.Y(_1928_),
    .A(_1926_),
    .B(_1927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5086_ (.B(_1928_),
    .A(_1925_),
    .X(_1929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5087_ (.A(_1908_),
    .B_N(_1929_),
    .Y(_1930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5088_ (.B(_1929_),
    .A(_1908_),
    .X(_1931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5089_ (.A(_1924_),
    .B(_1931_),
    .Y(_1932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5090_ (.B(_1931_),
    .A(_1924_),
    .X(_1933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5091_ (.Y(_1934_),
    .A(_1911_),
    .B(_1933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5092_ (.Y(_1935_),
    .A(_1911_),
    .B(_1933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5093_ (.B(_1935_),
    .A(_1923_),
    .X(_1936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5094_ (.A(_1922_),
    .B(_1936_),
    .X(_1937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5095_ (.Y(_1938_),
    .A(_1922_),
    .B(_1936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5096_ (.A(_1938_),
    .B_N(_1921_),
    .Y(_1939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5097_ (.B(_1938_),
    .A(_1921_),
    .X(_1940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5098_ (.B1(net475),
    .VDD(VPWR),
    .Y(_1941_),
    .VSS(VGND),
    .A1(net585),
    .A2(net864));
 sg13g2_a21oi_1 _5099_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net585),
    .A2(_1940_),
    .Y(_0275_),
    .B1(_1941_));
 sg13g2_nand2_1 _5100_ (.Y(_1942_),
    .A(\mydesign.pe_weights[33] ),
    .B(\mydesign.pe_inputs[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5101_ (.B1(_1926_),
    .VDD(VPWR),
    .Y(_1943_),
    .VSS(VGND),
    .A1(_1925_),
    .A2(_1928_));
 sg13g2_nand2_1 _5102_ (.Y(_1944_),
    .A(\mydesign.pe_weights[35] ),
    .B(\mydesign.pe_inputs[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5103_ (.B(net530),
    .C(\mydesign.pe_inputs[22] ),
    .A(\mydesign.accum[36] ),
    .Y(_1945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5104_ (.A2(\mydesign.pe_inputs[22] ),
    .A1(net530),
    .B1(\mydesign.accum[36] ),
    .X(_1946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5105_ (.Y(_1947_),
    .A(_1945_),
    .B(_1946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5106_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1948_),
    .B(_1947_),
    .A(_1944_));
 sg13g2_xor2_1 _5107_ (.B(_1947_),
    .A(_1944_),
    .X(_1949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5108_ (.Y(_1950_),
    .A(_1943_),
    .B(_1949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5109_ (.Y(_1951_),
    .A(_1943_),
    .B(_1949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5110_ (.B(_1951_),
    .A(_1942_),
    .X(_1952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5111_ (.B1(_1952_),
    .VDD(VPWR),
    .Y(_1953_),
    .VSS(VGND),
    .A1(_1930_),
    .A2(_1932_));
 sg13g2_or3_1 _5112_ (.A(_1930_),
    .B(_1932_),
    .C(_1952_),
    .X(_1954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5113_ (.A(_1953_),
    .B(_1954_),
    .X(_1955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5114_ (.B1(_1934_),
    .VDD(VPWR),
    .Y(_1956_),
    .VSS(VGND),
    .A1(_1923_),
    .A2(_1935_));
 sg13g2_nand2_1 _5115_ (.Y(_1957_),
    .A(_1955_),
    .B(_1956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5116_ (.B(_1956_),
    .A(_1955_),
    .X(_1958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5117_ (.A(_1937_),
    .B(_1939_),
    .C(_1958_),
    .X(_1959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5118_ (.B1(_1958_),
    .VDD(VPWR),
    .Y(_1960_),
    .VSS(VGND),
    .A1(_1937_),
    .A2(_1939_));
 sg13g2_a21oi_1 _5119_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1959_),
    .A2(_1960_),
    .Y(_1961_),
    .B1(net503));
 sg13g2_o21ai_1 _5120_ (.B1(net475),
    .VDD(VPWR),
    .Y(_1962_),
    .VSS(VGND),
    .A1(net584),
    .A2(net1002));
 sg13g2_nor2_1 _5121_ (.A(_1961_),
    .B(_1962_),
    .Y(_0276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5122_ (.B1(_1950_),
    .VDD(VPWR),
    .Y(_1963_),
    .VSS(VGND),
    .A1(_1942_),
    .A2(_1951_));
 sg13g2_nand2_1 _5123_ (.Y(_1964_),
    .A(\mydesign.pe_weights[35] ),
    .B(\mydesign.pe_inputs[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5124_ (.B(net530),
    .C(\mydesign.pe_inputs[23] ),
    .A(\mydesign.accum[37] ),
    .Y(_1965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5125_ (.A2(\mydesign.pe_inputs[23] ),
    .A1(net530),
    .B1(\mydesign.accum[37] ),
    .X(_1966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5126_ (.Y(_1967_),
    .A(_1965_),
    .B(_1966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5127_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1968_),
    .B(_1967_),
    .A(_1964_));
 sg13g2_xnor2_1 _5128_ (.Y(_1969_),
    .A(_1964_),
    .B(_1967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5129_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1945_),
    .A2(_1948_),
    .Y(_1970_),
    .B1(_1969_));
 sg13g2_nand3_1 _5130_ (.B(_1948_),
    .C(_1969_),
    .A(_1945_),
    .Y(_1971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5131_ (.A(_1970_),
    .B_N(_1971_),
    .Y(_1972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5132_ (.Y(_1973_),
    .A(_1963_),
    .B(_1972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5133_ (.Y(_1974_),
    .A(_1963_),
    .B(_1972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5134_ (.A(_1953_),
    .B(_1974_),
    .Y(_1975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5135_ (.Y(_1976_),
    .A(_1953_),
    .B(_1974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5136_ (.X(_1977_),
    .A(_1957_),
    .B(_1960_),
    .C(_1976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _5137_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1976_),
    .Y(_1978_),
    .A2(_1960_),
    .A1(_1957_));
 sg13g2_o21ai_1 _5138_ (.B1(net584),
    .VDD(VPWR),
    .Y(_1979_),
    .VSS(VGND),
    .A1(_1977_),
    .A2(_1978_));
 sg13g2_o21ai_1 _5139_ (.B1(net475),
    .VDD(VPWR),
    .Y(_1980_),
    .VSS(VGND),
    .A1(net584),
    .A2(net1005));
 sg13g2_nor2b_1 _5140_ (.A(_1980_),
    .B_N(_1979_),
    .Y(_0277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5141_ (.B(\mydesign.pe_weights[35] ),
    .C(\mydesign.pe_inputs[23] ),
    .A(\mydesign.accum[38] ),
    .Y(_1981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5142_ (.A2(\mydesign.pe_inputs[23] ),
    .A1(\mydesign.pe_weights[35] ),
    .B1(\mydesign.accum[38] ),
    .X(_1982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5143_ (.Y(_1983_),
    .A(_1981_),
    .B(_1982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5144_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1965_),
    .A2(_1968_),
    .Y(_1984_),
    .B1(_1983_));
 sg13g2_nand3_1 _5145_ (.B(_1968_),
    .C(_1983_),
    .A(_1965_),
    .Y(_1985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5146_ (.Y(_1986_),
    .B(_1985_),
    .A_N(_1984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5147_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1963_),
    .A2(_1971_),
    .Y(_1987_),
    .B1(_1970_));
 sg13g2_xor2_1 _5148_ (.B(_1987_),
    .A(_1986_),
    .X(_1988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5149_ (.A(_1975_),
    .B(_1978_),
    .C(_1988_),
    .Y(_1989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5150_ (.B1(_1988_),
    .VDD(VPWR),
    .Y(_1990_),
    .VSS(VGND),
    .A1(_1975_),
    .A2(_1978_));
 sg13g2_nand2b_1 _5151_ (.Y(_1991_),
    .B(_1990_),
    .A_N(_1989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5152_ (.B1(net474),
    .VDD(VPWR),
    .Y(_1992_),
    .VSS(VGND),
    .A1(net575),
    .A2(net826));
 sg13g2_a21oi_1 _5153_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net575),
    .A2(_1991_),
    .Y(_0278_),
    .B1(_1992_));
 sg13g2_o21ai_1 _5154_ (.B1(_1990_),
    .VDD(VPWR),
    .Y(_1993_),
    .VSS(VGND),
    .A1(_1973_),
    .A2(_1986_));
 sg13g2_a21oi_1 _5155_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1970_),
    .A2(_1985_),
    .Y(_1994_),
    .B1(_1984_));
 sg13g2_xnor2_1 _5156_ (.Y(_1995_),
    .A(net889),
    .B(_1981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5157_ (.Y(_1996_),
    .A(_1994_),
    .B(_1995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5158_ (.Y(_1997_),
    .A(_1993_),
    .B(_1996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5159_ (.B1(net474),
    .VDD(VPWR),
    .Y(_1998_),
    .VSS(VGND),
    .A1(net575),
    .A2(net889));
 sg13g2_a21oi_1 _5160_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net575),
    .A2(_1997_),
    .Y(_0279_),
    .B1(_1998_));
 sg13g2_nor2b_1 _5161_ (.A(\mydesign.inputs[3][4] ),
    .B_N(net549),
    .Y(_1999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5162_ (.A(net549),
    .B(\mydesign.inputs[3][8] ),
    .Y(_2000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5163_ (.A(_0397_),
    .B(_1999_),
    .C(_2000_),
    .Y(_2001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5164_ (.X(_2002_),
    .A(net549),
    .B(\mydesign.inputs[3][12] ),
    .C(_0392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5165_ (.X(_2003_),
    .A(net541),
    .B(\mydesign.inputs[3][0] ),
    .C(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5166_ (.A(_2001_),
    .B(_2002_),
    .C(_2003_),
    .X(_2004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5167_ (.B1(net625),
    .VDD(VPWR),
    .Y(_2005_),
    .VSS(VGND),
    .A1(net489),
    .A2(_2004_));
 sg13g2_a21oi_1 _5168_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2527_),
    .A2(net494),
    .Y(_0280_),
    .B1(_2005_));
 sg13g2_nand2b_1 _5169_ (.Y(_2006_),
    .B(\mydesign.inputs[3][9] ),
    .A_N(net549),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5170_ (.Y(_2007_),
    .A(net549),
    .B(\mydesign.inputs[3][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5171_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2006_),
    .A2(_2007_),
    .Y(_2008_),
    .B1(_0397_));
 sg13g2_a221oi_1 _5172_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\mydesign.inputs[3][13] ),
    .C1(_2008_),
    .B1(_0395_),
    .A1(\mydesign.inputs[3][1] ),
    .Y(_2009_),
    .A2(net454));
 sg13g2_inv_1 _5173_ (.VDD(VPWR),
    .Y(_2010_),
    .A(_2009_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5174_ (.B1(net634),
    .VDD(VPWR),
    .Y(_2011_),
    .VSS(VGND),
    .A1(net976),
    .A2(net445));
 sg13g2_a21oi_1 _5175_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net445),
    .A2(_2009_),
    .Y(_0281_),
    .B1(_2011_));
 sg13g2_nor2_1 _5176_ (.A(net497),
    .B(\mydesign.inputs[3][6] ),
    .Y(_2012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5177_ (.B1(net459),
    .VDD(VPWR),
    .Y(_2013_),
    .VSS(VGND),
    .A1(net549),
    .A2(\mydesign.inputs[3][10] ));
 sg13g2_a22oi_1 _5178_ (.Y(_2014_),
    .B1(_0395_),
    .B2(\mydesign.inputs[3][14] ),
    .A2(net454),
    .A1(\mydesign.inputs[3][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5179_ (.B1(_2014_),
    .VDD(VPWR),
    .Y(_2015_),
    .VSS(VGND),
    .A1(_2012_),
    .A2(_2013_));
 sg13g2_o21ai_1 _5180_ (.B1(net625),
    .VDD(VPWR),
    .Y(_2016_),
    .VSS(VGND),
    .A1(net487),
    .A2(_2015_));
 sg13g2_a21oi_1 _5181_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2526_),
    .A2(net494),
    .Y(_0282_),
    .B1(_2016_));
 sg13g2_nor2_1 _5182_ (.A(net497),
    .B(\mydesign.inputs[3][7] ),
    .Y(_2017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5183_ (.B1(net459),
    .VDD(VPWR),
    .Y(_2018_),
    .VSS(VGND),
    .A1(net549),
    .A2(\mydesign.inputs[3][11] ));
 sg13g2_a22oi_1 _5184_ (.Y(_2019_),
    .B1(_0395_),
    .B2(\mydesign.inputs[3][15] ),
    .A2(_2596_),
    .A1(\mydesign.inputs[3][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5185_ (.B1(_2019_),
    .VDD(VPWR),
    .Y(_2020_),
    .VSS(VGND),
    .A1(_2017_),
    .A2(_2018_));
 sg13g2_o21ai_1 _5186_ (.B1(net625),
    .VDD(VPWR),
    .Y(_2021_),
    .VSS(VGND),
    .A1(net487),
    .A2(_2020_));
 sg13g2_a21oi_1 _5187_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2525_),
    .A2(net494),
    .Y(_0283_),
    .B1(_2021_));
 sg13g2_and2_1 _5188_ (.A(net891),
    .B(_2004_),
    .X(_2022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5189_ (.Y(_2023_),
    .A(net563),
    .B(_2022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5190_ (.B(_2023_),
    .A(net979),
    .X(_2024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5191_ (.A(net462),
    .B(_2024_),
    .Y(_0284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5192_ (.B(\mydesign.pe_weights[29] ),
    .C(_2004_),
    .A(\mydesign.accum[25] ),
    .Y(_2025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5193_ (.A2(_2004_),
    .A1(\mydesign.pe_weights[29] ),
    .B1(\mydesign.accum[25] ),
    .X(_2026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5194_ (.Y(_2027_),
    .A(_2025_),
    .B(_2026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5195_ (.Y(_2028_),
    .A(net891),
    .B(_2010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5196_ (.A(_2027_),
    .B(_2028_),
    .Y(_2029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5197_ (.B(_2028_),
    .A(_2027_),
    .X(_2030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _5198_ (.X(_2031_),
    .A(\mydesign.accum[24] ),
    .B(_2022_),
    .C(_2030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5199_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[24] ),
    .A2(_2022_),
    .Y(_2032_),
    .B1(_2030_));
 sg13g2_or2_1 _5200_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2033_),
    .B(_2032_),
    .A(_2031_));
 sg13g2_o21ai_1 _5201_ (.B1(net466),
    .VDD(VPWR),
    .Y(_2034_),
    .VSS(VGND),
    .A1(net563),
    .A2(net954));
 sg13g2_a21oi_1 _5202_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net563),
    .A2(_2033_),
    .Y(_0285_),
    .B1(_2034_));
 sg13g2_nand2_1 _5203_ (.Y(_2035_),
    .A(\mydesign.pe_weights[28] ),
    .B(_2015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5204_ (.X(_2036_),
    .A(\mydesign.accum[26] ),
    .B(\mydesign.pe_weights[30] ),
    .C(_2004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5205_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[30] ),
    .A2(_2004_),
    .Y(_2037_),
    .B1(\mydesign.accum[26] ));
 sg13g2_or2_1 _5206_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2038_),
    .B(_2037_),
    .A(_2036_));
 sg13g2_nand2_1 _5207_ (.Y(_2039_),
    .A(\mydesign.pe_weights[29] ),
    .B(_2010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5208_ (.A(_2038_),
    .B(_2039_),
    .Y(_2040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5209_ (.B(_2039_),
    .A(_2038_),
    .X(_2041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5210_ (.Y(_2042_),
    .B(_2041_),
    .A_N(_2025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5211_ (.Y(_2043_),
    .A(_2025_),
    .B(_2041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5212_ (.Y(_2044_),
    .B(_2043_),
    .A_N(_2035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5213_ (.Y(_2045_),
    .A(_2035_),
    .B(_2043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5214_ (.A(_2029_),
    .B(_2045_),
    .X(_2046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5215_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2047_),
    .B(_2045_),
    .A(_2029_));
 sg13g2_nand2b_1 _5216_ (.Y(_2048_),
    .B(_2047_),
    .A_N(_2046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5217_ (.B(_2048_),
    .A(_2031_),
    .X(_2049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5218_ (.B1(net466),
    .VDD(VPWR),
    .Y(_2050_),
    .VSS(VGND),
    .A1(net563),
    .A2(net923));
 sg13g2_a21oi_1 _5219_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net563),
    .A2(_2049_),
    .Y(_0286_),
    .B1(_2050_));
 sg13g2_a21oi_1 _5220_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2031_),
    .A2(_2047_),
    .Y(_2051_),
    .B1(_2046_));
 sg13g2_nand2_1 _5221_ (.Y(_2052_),
    .A(_2042_),
    .B(_2044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5222_ (.Y(_2053_),
    .A(\mydesign.pe_weights[28] ),
    .B(_2020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5223_ (.VDD(VPWR),
    .Y(_2054_),
    .A(_2053_),
    .VSS(VGND));
 sg13g2_and2_1 _5224_ (.A(\mydesign.pe_weights[29] ),
    .B(_2015_),
    .X(_2055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5225_ (.A(_2009_),
    .B_N(\mydesign.pe_weights[30] ),
    .Y(_2056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5226_ (.B(\mydesign.pe_weights[31] ),
    .C(_2004_),
    .A(\mydesign.accum[27] ),
    .Y(_2057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5227_ (.A2(_2004_),
    .A1(\mydesign.pe_weights[31] ),
    .B1(\mydesign.accum[27] ),
    .X(_2058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5228_ (.B(_2057_),
    .C(_2058_),
    .A(_2056_),
    .Y(_2059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5229_ (.A2(_2058_),
    .A1(_2057_),
    .B1(_2056_),
    .X(_2060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5230_ (.B(_2059_),
    .C(_2060_),
    .A(_2036_),
    .Y(_2061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5231_ (.A2(_2060_),
    .A1(_2059_),
    .B1(_2036_),
    .X(_2062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5232_ (.B(_2061_),
    .C(_2062_),
    .A(_2055_),
    .Y(_2063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5233_ (.A2(_2062_),
    .A1(_2061_),
    .B1(_2055_),
    .X(_2064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5234_ (.B(_2063_),
    .C(_2064_),
    .A(_2040_),
    .Y(_2065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5235_ (.A2(_2064_),
    .A1(_2063_),
    .B1(_2040_),
    .X(_2066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5236_ (.B(_2065_),
    .C(_2066_),
    .A(_2054_),
    .Y(_2067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5237_ (.A2(_2066_),
    .A1(_2065_),
    .B1(_2054_),
    .X(_2068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5238_ (.Y(_2069_),
    .A(_2067_),
    .B(_2068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5239_ (.B(_2067_),
    .C(_2068_),
    .A(_2052_),
    .Y(_2070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5240_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2067_),
    .A2(_2068_),
    .Y(_2071_),
    .B1(_2052_));
 sg13g2_xnor2_1 _5241_ (.Y(_2072_),
    .A(_2052_),
    .B(_2069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5242_ (.Y(_2073_),
    .A(_2051_),
    .B(_2072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5243_ (.B1(net466),
    .VDD(VPWR),
    .Y(_2074_),
    .VSS(VGND),
    .A1(net499),
    .A2(_2073_));
 sg13g2_a21oi_1 _5244_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net499),
    .A2(_2528_),
    .Y(_0287_),
    .B1(_2074_));
 sg13g2_o21ai_1 _5245_ (.B1(_2070_),
    .VDD(VPWR),
    .Y(_2075_),
    .VSS(VGND),
    .A1(_2051_),
    .A2(_2071_));
 sg13g2_nand2_1 _5246_ (.Y(_2076_),
    .A(_2065_),
    .B(_2067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5247_ (.Y(_2077_),
    .A(_2061_),
    .B(_2063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5248_ (.Y(_2078_),
    .A(\mydesign.pe_weights[29] ),
    .B(_2020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5249_ (.Y(_2079_),
    .A(_2057_),
    .B(_2059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5250_ (.Y(_2080_),
    .A(\mydesign.pe_weights[30] ),
    .B(_2015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5251_ (.A(_2009_),
    .B_N(\mydesign.pe_weights[31] ),
    .Y(_2081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5252_ (.Y(_2082_),
    .A(\mydesign.accum[28] ),
    .B(_2081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5253_ (.A(_2080_),
    .B(_2082_),
    .Y(_2083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5254_ (.B(_2082_),
    .A(_2080_),
    .X(_2084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5255_ (.Y(_2085_),
    .A(_2079_),
    .B(_2084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5256_ (.Y(_2086_),
    .A(_2079_),
    .B(_2084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5257_ (.B(_2086_),
    .A(_2078_),
    .X(_2087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5258_ (.Y(_2088_),
    .A(_2077_),
    .B(_2087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5259_ (.Y(_2089_),
    .A(_2077_),
    .B(_2087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5260_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2065_),
    .A2(_2067_),
    .Y(_2090_),
    .B1(_2089_));
 sg13g2_xnor2_1 _5261_ (.Y(_2091_),
    .A(_2076_),
    .B(_2089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5262_ (.Y(_2092_),
    .A(_2075_),
    .B(_2091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5263_ (.B1(net464),
    .VDD(VPWR),
    .Y(_2093_),
    .VSS(VGND),
    .A1(net565),
    .A2(net1012));
 sg13g2_a21oi_1 _5264_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net565),
    .A2(_2092_),
    .Y(_0288_),
    .B1(_2093_));
 sg13g2_a21oi_1 _5265_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2075_),
    .A2(_2091_),
    .Y(_2094_),
    .B1(_2090_));
 sg13g2_o21ai_1 _5266_ (.B1(_2085_),
    .VDD(VPWR),
    .Y(_2095_),
    .VSS(VGND),
    .A1(_2078_),
    .A2(_2086_));
 sg13g2_nand2_1 _5267_ (.Y(_2096_),
    .A(\mydesign.pe_weights[30] ),
    .B(_2020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5268_ (.B(\mydesign.pe_weights[31] ),
    .C(_2015_),
    .A(\mydesign.accum[29] ),
    .Y(_2097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5269_ (.A2(_2015_),
    .A1(\mydesign.pe_weights[31] ),
    .B1(\mydesign.accum[29] ),
    .X(_2098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5270_ (.Y(_2099_),
    .A(_2097_),
    .B(_2098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5271_ (.B(_2099_),
    .A(_2096_),
    .X(_2100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5272_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[28] ),
    .A2(_2081_),
    .Y(_2101_),
    .B1(_2083_));
 sg13g2_nand2b_1 _5273_ (.Y(_2102_),
    .B(_2100_),
    .A_N(_2101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5274_ (.Y(_2103_),
    .A(_2100_),
    .B(_2101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5275_ (.Y(_2104_),
    .A(_2095_),
    .B(_2103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5276_ (.Y(_2105_),
    .A(_2095_),
    .B(_2103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5277_ (.A(_2088_),
    .B(_2105_),
    .X(_2106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5278_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2107_),
    .B(_2105_),
    .A(_2088_));
 sg13g2_nand2b_1 _5279_ (.Y(_2108_),
    .B(_2107_),
    .A_N(_2106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5280_ (.Y(_2109_),
    .A(_2094_),
    .B(_2108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5281_ (.B1(net465),
    .VDD(VPWR),
    .Y(_2110_),
    .VSS(VGND),
    .A1(net565),
    .A2(net890));
 sg13g2_a21oi_1 _5282_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net565),
    .A2(_2109_),
    .Y(_0289_),
    .B1(_2110_));
 sg13g2_a21oi_1 _5283_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_weights[31] ),
    .A2(_2020_),
    .Y(_2111_),
    .B1(\mydesign.accum[30] ));
 sg13g2_nand3_1 _5284_ (.B(\mydesign.pe_weights[31] ),
    .C(_2020_),
    .A(\mydesign.accum[30] ),
    .Y(_2112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5285_ (.Y(_2113_),
    .B(_2112_),
    .A_N(_2111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5286_ (.B1(_2097_),
    .VDD(VPWR),
    .Y(_2114_),
    .VSS(VGND),
    .A1(_2096_),
    .A2(_2099_));
 sg13g2_inv_1 _5287_ (.VDD(VPWR),
    .Y(_2115_),
    .A(_2114_),
    .VSS(VGND));
 sg13g2_xnor2_1 _5288_ (.Y(_2116_),
    .A(_2113_),
    .B(_2114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5289_ (.Y(_2117_),
    .B(_2116_),
    .A_N(_2102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5290_ (.Y(_2118_),
    .A(_2102_),
    .B(_2116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5291_ (.A(_2104_),
    .B_N(_2118_),
    .Y(_2119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5292_ (.Y(_2120_),
    .A(_2104_),
    .B(_2118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5293_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2094_),
    .A2(_2107_),
    .Y(_2121_),
    .B1(_2106_));
 sg13g2_xnor2_1 _5294_ (.Y(_2122_),
    .A(_2120_),
    .B(_2121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5295_ (.B1(net470),
    .VDD(VPWR),
    .Y(_2123_),
    .VSS(VGND),
    .A1(net568),
    .A2(net945));
 sg13g2_a21oi_1 _5296_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net568),
    .A2(_2122_),
    .Y(_0290_),
    .B1(_2123_));
 sg13g2_a21oi_1 _5297_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2120_),
    .A2(_2121_),
    .Y(_2124_),
    .B1(_2119_));
 sg13g2_o21ai_1 _5298_ (.B1(_2112_),
    .VDD(VPWR),
    .Y(_2125_),
    .VSS(VGND),
    .A1(_2111_),
    .A2(_2115_));
 sg13g2_xor2_1 _5299_ (.B(_2125_),
    .A(net837),
    .X(_2126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5300_ (.Y(_2127_),
    .A(_2117_),
    .B(_2126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5301_ (.B(_2127_),
    .A(_2124_),
    .X(_2128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5302_ (.B1(net470),
    .VDD(VPWR),
    .Y(_2129_),
    .VSS(VGND),
    .A1(net568),
    .A2(net837));
 sg13g2_a21oi_1 _5303_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net567),
    .A2(_2128_),
    .Y(_0291_),
    .B1(_2129_));
 sg13g2_nand2_2 _5304_ (.Y(_2130_),
    .A(net611),
    .B(_2640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5305_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net611),
    .A2(_2640_),
    .Y(_2131_),
    .B1(net608));
 sg13g2_nand2_1 _5306_ (.Y(_2132_),
    .A(net695),
    .B(_2131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5307_ (.B1(_2132_),
    .VDD(VPWR),
    .Y(_0292_),
    .VSS(VGND),
    .A1(net603),
    .A2(_2130_));
 sg13g2_nand2_1 _5308_ (.Y(_2133_),
    .A(net660),
    .B(_2131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5309_ (.B1(_2133_),
    .VDD(VPWR),
    .Y(_0293_),
    .VSS(VGND),
    .A1(net601),
    .A2(_2130_));
 sg13g2_nand2_1 _5310_ (.Y(_2134_),
    .A(net427),
    .B(_2131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5311_ (.B1(_2134_),
    .VDD(VPWR),
    .Y(_0294_),
    .VSS(VGND),
    .A1(net599),
    .A2(_2130_));
 sg13g2_nand2_1 _5312_ (.Y(_2135_),
    .A(net656),
    .B(_2131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5313_ (.B1(_2135_),
    .VDD(VPWR),
    .Y(_0295_),
    .VSS(VGND),
    .A1(net597),
    .A2(_2130_));
 sg13g2_o21ai_1 _5314_ (.B1(net638),
    .VDD(VPWR),
    .Y(_2136_),
    .VSS(VGND),
    .A1(net521),
    .A2(net450));
 sg13g2_a21oi_1 _5315_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2527_),
    .A2(net449),
    .Y(_0296_),
    .B1(_2136_));
 sg13g2_o21ai_1 _5316_ (.B1(net634),
    .VDD(VPWR),
    .Y(_2137_),
    .VSS(VGND),
    .A1(net976),
    .A2(net493));
 sg13g2_a21oi_1 _5317_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2523_),
    .A2(net493),
    .Y(_0297_),
    .B1(_2137_));
 sg13g2_o21ai_1 _5318_ (.B1(net638),
    .VDD(VPWR),
    .Y(_2138_),
    .VSS(VGND),
    .A1(net832),
    .A2(net449));
 sg13g2_a21oi_1 _5319_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2526_),
    .A2(net449),
    .Y(_0298_),
    .B1(_2138_));
 sg13g2_o21ai_1 _5320_ (.B1(net638),
    .VDD(VPWR),
    .Y(_2139_),
    .VSS(VGND),
    .A1(net520),
    .A2(net450));
 sg13g2_a21oi_1 _5321_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2525_),
    .A2(net449),
    .Y(_0299_),
    .B1(_2139_));
 sg13g2_and3_1 _5322_ (.X(_2140_),
    .A(net591),
    .B(net522),
    .C(\mydesign.pe_weights[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5323_ (.B1(net481),
    .VDD(VPWR),
    .Y(_2141_),
    .VSS(VGND),
    .A1(net758),
    .A2(_2140_));
 sg13g2_a21oi_1 _5324_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net758),
    .A2(_2140_),
    .Y(_0300_),
    .B1(_2141_));
 sg13g2_and3_2 _5325_ (.X(_2142_),
    .A(\mydesign.accum[17] ),
    .B(net522),
    .C(\mydesign.pe_weights[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5326_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net522),
    .A2(\mydesign.pe_weights[25] ),
    .Y(_2143_),
    .B1(\mydesign.accum[17] ));
 sg13g2_nand2_1 _5327_ (.Y(_2144_),
    .A(\mydesign.pe_inputs[13] ),
    .B(\mydesign.pe_weights[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5328_ (.A(_2142_),
    .B(_2143_),
    .C(_2144_),
    .Y(_2145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5329_ (.B1(_2144_),
    .VDD(VPWR),
    .Y(_2146_),
    .VSS(VGND),
    .A1(_2142_),
    .A2(_2143_));
 sg13g2_nor2b_1 _5330_ (.A(_2145_),
    .B_N(_2146_),
    .Y(_2147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5331_ (.B(net522),
    .C(\mydesign.pe_weights[24] ),
    .A(net758),
    .Y(_2148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5332_ (.B(net522),
    .C(\mydesign.pe_weights[24] ),
    .A(net758),
    .Y(_2149_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2147_));
 sg13g2_xor2_1 _5333_ (.B(_2148_),
    .A(_2147_),
    .X(_2150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5334_ (.B1(net481),
    .VDD(VPWR),
    .Y(_2151_),
    .VSS(VGND),
    .A1(net591),
    .A2(net1029));
 sg13g2_a21oi_1 _5335_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net591),
    .A2(_2150_),
    .Y(_0301_),
    .B1(_2151_));
 sg13g2_nand2_1 _5336_ (.Y(_2152_),
    .A(\mydesign.pe_inputs[14] ),
    .B(\mydesign.pe_weights[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5337_ (.Y(_2153_),
    .A(\mydesign.pe_inputs[13] ),
    .B(\mydesign.pe_weights[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5338_ (.B(net522),
    .C(\mydesign.pe_weights[26] ),
    .A(\mydesign.accum[18] ),
    .Y(_2154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5339_ (.A2(\mydesign.pe_weights[26] ),
    .A1(net522),
    .B1(\mydesign.accum[18] ),
    .X(_2155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5340_ (.Y(_2156_),
    .A(_2154_),
    .B(_2155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5341_ (.A(_2153_),
    .B(_2156_),
    .Y(_2157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5342_ (.B(_2156_),
    .A(_2153_),
    .X(_2158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5343_ (.Y(_2159_),
    .A(_2142_),
    .B(_2158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5344_ (.A(_2142_),
    .B(_2158_),
    .Y(_2160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5345_ (.B(_2158_),
    .A(_2142_),
    .X(_2161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5346_ (.Y(_2162_),
    .A(_2152_),
    .B(_2161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5347_ (.Y(_2163_),
    .A(_2145_),
    .B(_2162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5348_ (.Y(_2164_),
    .A(_2145_),
    .B(_2162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5349_ (.Y(_2165_),
    .A(_2149_),
    .B(_2164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5350_ (.B1(net481),
    .VDD(VPWR),
    .Y(_2166_),
    .VSS(VGND),
    .A1(net590),
    .A2(net1020));
 sg13g2_a21oi_1 _5351_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net591),
    .A2(_2165_),
    .Y(_0302_),
    .B1(_2166_));
 sg13g2_o21ai_1 _5352_ (.B1(_2163_),
    .VDD(VPWR),
    .Y(_2167_),
    .VSS(VGND),
    .A1(_2149_),
    .A2(_2164_));
 sg13g2_o21ai_1 _5353_ (.B1(_2159_),
    .VDD(VPWR),
    .Y(_2168_),
    .VSS(VGND),
    .A1(_2152_),
    .A2(_2160_));
 sg13g2_nand2_1 _5354_ (.Y(_2169_),
    .A(\mydesign.pe_inputs[15] ),
    .B(\mydesign.pe_weights[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5355_ (.Y(_2170_),
    .A(\mydesign.pe_inputs[14] ),
    .B(\mydesign.pe_weights[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5356_ (.Y(_2171_),
    .A(\mydesign.pe_inputs[13] ),
    .B(\mydesign.pe_weights[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5357_ (.B(\mydesign.pe_inputs[12] ),
    .C(net527),
    .A(\mydesign.accum[19] ),
    .Y(_2172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5358_ (.A2(net527),
    .A1(\mydesign.pe_inputs[12] ),
    .B1(\mydesign.accum[19] ),
    .X(_2173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5359_ (.Y(_2174_),
    .A(_2172_),
    .B(_2173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5360_ (.B(_2174_),
    .A(_2171_),
    .X(_2175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5361_ (.A(_2154_),
    .B_N(_2175_),
    .Y(_2176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5362_ (.B(_2175_),
    .A(_2154_),
    .X(_2177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5363_ (.A(_2170_),
    .B(_2177_),
    .Y(_2178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5364_ (.B(_2177_),
    .A(_2170_),
    .X(_2179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5365_ (.Y(_2180_),
    .A(_2157_),
    .B(_2179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5366_ (.Y(_2181_),
    .A(_2157_),
    .B(_2179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5367_ (.B(_2181_),
    .A(_2169_),
    .X(_2182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5368_ (.A(_2168_),
    .B(_2182_),
    .X(_2183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5369_ (.Y(_2184_),
    .A(_2168_),
    .B(_2182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5370_ (.A(_2184_),
    .B_N(_2167_),
    .Y(_2185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5371_ (.B(_2184_),
    .A(_2167_),
    .X(_2186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5372_ (.B1(net481),
    .VDD(VPWR),
    .Y(_2187_),
    .VSS(VGND),
    .A1(net590),
    .A2(net992));
 sg13g2_a21oi_1 _5373_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net590),
    .A2(_2186_),
    .Y(_0303_),
    .B1(_2187_));
 sg13g2_nand2_1 _5374_ (.Y(_2188_),
    .A(\mydesign.pe_inputs[15] ),
    .B(\mydesign.pe_weights[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5375_ (.B1(_2172_),
    .VDD(VPWR),
    .Y(_2189_),
    .VSS(VGND),
    .A1(_2171_),
    .A2(_2174_));
 sg13g2_nand2_1 _5376_ (.Y(_2190_),
    .A(\mydesign.pe_inputs[14] ),
    .B(\mydesign.pe_weights[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5377_ (.B(\mydesign.pe_inputs[13] ),
    .C(net527),
    .A(\mydesign.accum[20] ),
    .Y(_2191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5378_ (.A2(net527),
    .A1(\mydesign.pe_inputs[13] ),
    .B1(\mydesign.accum[20] ),
    .X(_2192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5379_ (.Y(_2193_),
    .A(_2191_),
    .B(_2192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5380_ (.B(_2193_),
    .A(_2190_),
    .X(_2194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5381_ (.Y(_2195_),
    .A(_2189_),
    .B(_2194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5382_ (.Y(_2196_),
    .A(_2189_),
    .B(_2194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5383_ (.B(_2196_),
    .A(_2188_),
    .X(_2197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5384_ (.B1(_2197_),
    .VDD(VPWR),
    .Y(_2198_),
    .VSS(VGND),
    .A1(_2176_),
    .A2(_2178_));
 sg13g2_or3_1 _5385_ (.A(_2176_),
    .B(_2178_),
    .C(_2197_),
    .X(_2199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5386_ (.A(_2198_),
    .B(_2199_),
    .X(_2200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5387_ (.B1(_2180_),
    .VDD(VPWR),
    .Y(_2201_),
    .VSS(VGND),
    .A1(_2169_),
    .A2(_2181_));
 sg13g2_nand2_1 _5388_ (.Y(_2202_),
    .A(_2200_),
    .B(_2201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5389_ (.B(_2201_),
    .A(_2200_),
    .X(_2203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5390_ (.A(_2183_),
    .B(_2185_),
    .C(_2203_),
    .X(_2204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5391_ (.B1(_2203_),
    .VDD(VPWR),
    .Y(_2205_),
    .VSS(VGND),
    .A1(_2183_),
    .A2(_2185_));
 sg13g2_a21oi_1 _5392_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2204_),
    .A2(_2205_),
    .Y(_2206_),
    .B1(net503));
 sg13g2_o21ai_1 _5393_ (.B1(net481),
    .VDD(VPWR),
    .Y(_2207_),
    .VSS(VGND),
    .A1(net590),
    .A2(net1042));
 sg13g2_nor2_1 _5394_ (.A(_2206_),
    .B(_2207_),
    .Y(_0304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5395_ (.Y(_2208_),
    .A(\mydesign.pe_inputs[15] ),
    .B(\mydesign.pe_weights[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5396_ (.B(\mydesign.pe_inputs[14] ),
    .C(net527),
    .A(\mydesign.accum[21] ),
    .Y(_2209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5397_ (.A2(net527),
    .A1(\mydesign.pe_inputs[14] ),
    .B1(\mydesign.accum[21] ),
    .X(_2210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5398_ (.Y(_2211_),
    .A(_2209_),
    .B(_2210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5399_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2212_),
    .B(_2211_),
    .A(_2208_));
 sg13g2_xor2_1 _5400_ (.B(_2211_),
    .A(_2208_),
    .X(_2213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5401_ (.B1(_2191_),
    .VDD(VPWR),
    .Y(_2214_),
    .VSS(VGND),
    .A1(_2190_),
    .A2(_2193_));
 sg13g2_and2_1 _5402_ (.A(_2213_),
    .B(_2214_),
    .X(_2215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5403_ (.B(_2214_),
    .A(_2213_),
    .X(_2216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5404_ (.B1(_2195_),
    .VDD(VPWR),
    .Y(_2217_),
    .VSS(VGND),
    .A1(_2188_),
    .A2(_2196_));
 sg13g2_nand2_1 _5405_ (.Y(_2218_),
    .A(_2216_),
    .B(_2217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5406_ (.B(_2217_),
    .A(_2216_),
    .X(_2219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5407_ (.A(_2198_),
    .B_N(_2219_),
    .Y(_2220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5408_ (.B(_2219_),
    .A(_2198_),
    .X(_2221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5409_ (.X(_2222_),
    .A(_2202_),
    .B(_2205_),
    .C(_2221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5410_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2202_),
    .A2(_2205_),
    .Y(_2223_),
    .B1(_2221_));
 sg13g2_o21ai_1 _5411_ (.B1(net593),
    .VDD(VPWR),
    .Y(_2224_),
    .VSS(VGND),
    .A1(_2222_),
    .A2(_2223_));
 sg13g2_o21ai_1 _5412_ (.B1(net482),
    .VDD(VPWR),
    .Y(_2225_),
    .VSS(VGND),
    .A1(net590),
    .A2(net1035));
 sg13g2_nor2b_1 _5413_ (.A(_2225_),
    .B_N(_2224_),
    .Y(_0305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5414_ (.B(\mydesign.pe_inputs[15] ),
    .C(net527),
    .A(\mydesign.accum[22] ),
    .Y(_2226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5415_ (.A2(\mydesign.pe_weights[27] ),
    .A1(\mydesign.pe_inputs[15] ),
    .B1(\mydesign.accum[22] ),
    .X(_2227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5416_ (.Y(_2228_),
    .A(_2226_),
    .B(_2227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5417_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2209_),
    .A2(_2212_),
    .Y(_2229_),
    .B1(_2228_));
 sg13g2_nand3_1 _5418_ (.B(_2212_),
    .C(_2228_),
    .A(_2209_),
    .Y(_2230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5419_ (.Y(_2231_),
    .B(_2230_),
    .A_N(_2229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5420_ (.Y(_2232_),
    .B(_2218_),
    .A_N(_2215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5421_ (.Y(_2233_),
    .A(_2231_),
    .B(_2232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5422_ (.A(_2220_),
    .B(_2223_),
    .C(_2233_),
    .X(_2234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5423_ (.B1(_2233_),
    .VDD(VPWR),
    .Y(_2235_),
    .VSS(VGND),
    .A1(_2220_),
    .A2(_2223_));
 sg13g2_a21oi_1 _5424_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2234_),
    .A2(_2235_),
    .Y(_2236_),
    .B1(net502));
 sg13g2_o21ai_1 _5425_ (.B1(net482),
    .VDD(VPWR),
    .Y(_2237_),
    .VSS(VGND),
    .A1(net590),
    .A2(net915));
 sg13g2_nor2_1 _5426_ (.A(_2236_),
    .B(_2237_),
    .Y(_0306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5427_ (.B1(_2235_),
    .VDD(VPWR),
    .Y(_2238_),
    .VSS(VGND),
    .A1(_2218_),
    .A2(_2231_));
 sg13g2_a21oi_1 _5428_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2215_),
    .A2(_2230_),
    .Y(_2239_),
    .B1(_2229_));
 sg13g2_xnor2_1 _5429_ (.Y(_2240_),
    .A(net978),
    .B(_2226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5430_ (.Y(_2241_),
    .A(_2239_),
    .B(_2240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5431_ (.Y(_2242_),
    .A(_2238_),
    .B(_2241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5432_ (.B1(net482),
    .VDD(VPWR),
    .Y(_2243_),
    .VSS(VGND),
    .A1(net593),
    .A2(net978));
 sg13g2_a21oi_1 _5433_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net593),
    .A2(_2242_),
    .Y(_0307_),
    .B1(_2243_));
 sg13g2_o21ai_1 _5434_ (.B1(net635),
    .VDD(VPWR),
    .Y(_2244_),
    .VSS(VGND),
    .A1(net1065),
    .A2(net444));
 sg13g2_a21oi_1 _5435_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2524_),
    .A2(net444),
    .Y(_0308_),
    .B1(_2244_));
 sg13g2_o21ai_1 _5436_ (.B1(net635),
    .VDD(VPWR),
    .Y(_2245_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[5] ),
    .A2(net444));
 sg13g2_a21oi_1 _5437_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2523_),
    .A2(net444),
    .Y(_0309_),
    .B1(_2245_));
 sg13g2_o21ai_1 _5438_ (.B1(net635),
    .VDD(VPWR),
    .Y(_2246_),
    .VSS(VGND),
    .A1(\mydesign.pe_inputs[6] ),
    .A2(net444));
 sg13g2_a21oi_1 _5439_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2522_),
    .A2(net444),
    .Y(_0310_),
    .B1(_2246_));
 sg13g2_o21ai_1 _5440_ (.B1(net635),
    .VDD(VPWR),
    .Y(_2247_),
    .VSS(VGND),
    .A1(net946),
    .A2(net444));
 sg13g2_a21oi_1 _5441_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2521_),
    .A2(net445),
    .Y(_0311_),
    .B1(_2247_));
 sg13g2_and3_1 _5442_ (.X(_2248_),
    .A(net588),
    .B(net521),
    .C(\mydesign.pe_weights[20] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5443_ (.B1(net477),
    .VDD(VPWR),
    .Y(_2249_),
    .VSS(VGND),
    .A1(net729),
    .A2(_2248_));
 sg13g2_a21oi_1 _5444_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net729),
    .A2(_2248_),
    .Y(_0312_),
    .B1(_2249_));
 sg13g2_and3_2 _5445_ (.X(_2250_),
    .A(\mydesign.accum[9] ),
    .B(net521),
    .C(\mydesign.pe_weights[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5446_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net521),
    .A2(\mydesign.pe_weights[21] ),
    .Y(_2251_),
    .B1(\mydesign.accum[9] ));
 sg13g2_nand2_1 _5447_ (.Y(_2252_),
    .A(\mydesign.pe_inputs[9] ),
    .B(\mydesign.pe_weights[20] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5448_ (.A(_2250_),
    .B(_2251_),
    .C(_2252_),
    .Y(_2253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5449_ (.B1(_2252_),
    .VDD(VPWR),
    .Y(_2254_),
    .VSS(VGND),
    .A1(_2250_),
    .A2(_2251_));
 sg13g2_nor2b_1 _5450_ (.A(_2253_),
    .B_N(_2254_),
    .Y(_2255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5451_ (.B(net521),
    .C(\mydesign.pe_weights[20] ),
    .A(net729),
    .Y(_2256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5452_ (.B(net521),
    .C(\mydesign.pe_weights[20] ),
    .A(net729),
    .Y(_2257_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2255_));
 sg13g2_xor2_1 _5453_ (.B(_2256_),
    .A(_2255_),
    .X(_2258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5454_ (.B1(net477),
    .VDD(VPWR),
    .Y(_2259_),
    .VSS(VGND),
    .A1(net588),
    .A2(net928));
 sg13g2_a21oi_1 _5455_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net588),
    .A2(_2258_),
    .Y(_0313_),
    .B1(_2259_));
 sg13g2_nand2_1 _5456_ (.Y(_2260_),
    .A(\mydesign.pe_inputs[10] ),
    .B(\mydesign.pe_weights[20] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5457_ (.Y(_2261_),
    .A(\mydesign.pe_inputs[9] ),
    .B(\mydesign.pe_weights[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5458_ (.B(\mydesign.pe_inputs[8] ),
    .C(net525),
    .A(\mydesign.accum[10] ),
    .Y(_2262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5459_ (.A2(net525),
    .A1(\mydesign.pe_inputs[8] ),
    .B1(\mydesign.accum[10] ),
    .X(_2263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5460_ (.Y(_2264_),
    .A(_2262_),
    .B(_2263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5461_ (.A(_2261_),
    .B(_2264_),
    .Y(_2265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5462_ (.B(_2264_),
    .A(_2261_),
    .X(_2266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5463_ (.Y(_2267_),
    .A(_2250_),
    .B(_2266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5464_ (.A(_2250_),
    .B(_2266_),
    .Y(_2268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5465_ (.B(_2266_),
    .A(_2250_),
    .X(_2269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5466_ (.Y(_2270_),
    .A(_2260_),
    .B(_2269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5467_ (.Y(_2271_),
    .A(_2253_),
    .B(_2270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5468_ (.Y(_2272_),
    .A(_2253_),
    .B(_2270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5469_ (.Y(_2273_),
    .A(_2257_),
    .B(_2272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5470_ (.B1(net477),
    .VDD(VPWR),
    .Y(_2274_),
    .VSS(VGND),
    .A1(net588),
    .A2(net1038));
 sg13g2_a21oi_1 _5471_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net588),
    .A2(_2273_),
    .Y(_0314_),
    .B1(_2274_));
 sg13g2_o21ai_1 _5472_ (.B1(_2271_),
    .VDD(VPWR),
    .Y(_2275_),
    .VSS(VGND),
    .A1(_2257_),
    .A2(_2272_));
 sg13g2_o21ai_1 _5473_ (.B1(_2267_),
    .VDD(VPWR),
    .Y(_2276_),
    .VSS(VGND),
    .A1(_2260_),
    .A2(_2268_));
 sg13g2_nand2_1 _5474_ (.Y(_2277_),
    .A(net520),
    .B(\mydesign.pe_weights[20] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5475_ (.Y(_2278_),
    .A(\mydesign.pe_inputs[10] ),
    .B(\mydesign.pe_weights[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5476_ (.Y(_2279_),
    .A(net521),
    .B(\mydesign.pe_weights[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5477_ (.B(\mydesign.pe_inputs[9] ),
    .C(\mydesign.pe_weights[22] ),
    .A(\mydesign.accum[11] ),
    .Y(_2280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5478_ (.A2(\mydesign.pe_weights[22] ),
    .A1(\mydesign.pe_inputs[9] ),
    .B1(\mydesign.accum[11] ),
    .X(_2281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5479_ (.Y(_2282_),
    .A(_2280_),
    .B(_2281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5480_ (.B(_2282_),
    .A(_2279_),
    .X(_2283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5481_ (.A(_2262_),
    .B_N(_2283_),
    .Y(_2284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5482_ (.B(_2283_),
    .A(_2262_),
    .X(_2285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5483_ (.A(_2278_),
    .B(_2285_),
    .Y(_2286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5484_ (.B(_2285_),
    .A(_2278_),
    .X(_2287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5485_ (.Y(_2288_),
    .A(_2265_),
    .B(_2287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5486_ (.Y(_2289_),
    .A(_2265_),
    .B(_2287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5487_ (.B(_2289_),
    .A(_2277_),
    .X(_2290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5488_ (.A(_2276_),
    .B(_2290_),
    .X(_2291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5489_ (.Y(_2292_),
    .A(_2276_),
    .B(_2290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5490_ (.A(_2292_),
    .B_N(_2275_),
    .Y(_2293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5491_ (.B(_2292_),
    .A(_2275_),
    .X(_2294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5492_ (.B1(net478),
    .VDD(VPWR),
    .Y(_2295_),
    .VSS(VGND),
    .A1(net588),
    .A2(net970));
 sg13g2_a21oi_1 _5493_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net588),
    .A2(_2294_),
    .Y(_0315_),
    .B1(_2295_));
 sg13g2_nand2_1 _5494_ (.Y(_2296_),
    .A(net520),
    .B(\mydesign.pe_weights[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5495_ (.B1(_2280_),
    .VDD(VPWR),
    .Y(_2297_),
    .VSS(VGND),
    .A1(_2279_),
    .A2(_2282_));
 sg13g2_nand2_1 _5496_ (.Y(_2298_),
    .A(\mydesign.pe_inputs[9] ),
    .B(\mydesign.pe_weights[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5497_ (.B(\mydesign.pe_inputs[10] ),
    .C(net525),
    .A(\mydesign.accum[12] ),
    .Y(_2299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5498_ (.A2(net525),
    .A1(\mydesign.pe_inputs[10] ),
    .B1(\mydesign.accum[12] ),
    .X(_2300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5499_ (.Y(_2301_),
    .A(_2299_),
    .B(_2300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5500_ (.B(_2301_),
    .A(_2298_),
    .X(_2302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5501_ (.Y(_2303_),
    .A(_2297_),
    .B(_2302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5502_ (.Y(_2304_),
    .A(_2297_),
    .B(_2302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5503_ (.B(_2304_),
    .A(_2296_),
    .X(_2305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5504_ (.B1(_2305_),
    .VDD(VPWR),
    .Y(_2306_),
    .VSS(VGND),
    .A1(_2284_),
    .A2(_2286_));
 sg13g2_or3_1 _5505_ (.A(_2284_),
    .B(_2286_),
    .C(_2305_),
    .X(_2307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5506_ (.A(_2306_),
    .B(_2307_),
    .X(_2308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5507_ (.B1(_2288_),
    .VDD(VPWR),
    .Y(_2309_),
    .VSS(VGND),
    .A1(_2277_),
    .A2(_2289_));
 sg13g2_nand2_1 _5508_ (.Y(_2310_),
    .A(_2308_),
    .B(_2309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5509_ (.B(_2309_),
    .A(_2308_),
    .X(_2311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5510_ (.A(_2291_),
    .B(_2293_),
    .C(_2311_),
    .Y(_2312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5511_ (.B1(_2311_),
    .VDD(VPWR),
    .Y(_2313_),
    .VSS(VGND),
    .A1(_2291_),
    .A2(_2293_));
 sg13g2_nand2b_1 _5512_ (.Y(_2314_),
    .B(_2313_),
    .A_N(_2312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5513_ (.B1(net481),
    .VDD(VPWR),
    .Y(_2315_),
    .VSS(VGND),
    .A1(net592),
    .A2(net1048));
 sg13g2_a21oi_1 _5514_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net592),
    .A2(_2314_),
    .Y(_0316_),
    .B1(_2315_));
 sg13g2_nand2_1 _5515_ (.Y(_2316_),
    .A(\mydesign.pe_inputs[10] ),
    .B(\mydesign.pe_weights[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5516_ (.X(_2317_),
    .A(\mydesign.accum[13] ),
    .B(net520),
    .C(net525),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5517_ (.B(net520),
    .C(net525),
    .A(\mydesign.accum[13] ),
    .Y(_2318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5518_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_inputs[11] ),
    .A2(net525),
    .Y(_2319_),
    .B1(\mydesign.accum[13] ));
 sg13g2_nor2_1 _5519_ (.A(_2317_),
    .B(_2319_),
    .Y(_2320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5520_ (.Y(_2321_),
    .A(_2316_),
    .B(_2320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5521_ (.B1(_2299_),
    .VDD(VPWR),
    .Y(_2322_),
    .VSS(VGND),
    .A1(_2298_),
    .A2(_2301_));
 sg13g2_xor2_1 _5522_ (.B(_2322_),
    .A(_2321_),
    .X(_2323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5523_ (.B1(_2303_),
    .VDD(VPWR),
    .Y(_2324_),
    .VSS(VGND),
    .A1(_2296_),
    .A2(_2304_));
 sg13g2_nand2_1 _5524_ (.Y(_2325_),
    .A(_2323_),
    .B(_2324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5525_ (.B(_2324_),
    .A(_2323_),
    .X(_2326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5526_ (.A(_2306_),
    .B_N(_2326_),
    .Y(_2327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5527_ (.B(_2326_),
    .A(_2306_),
    .X(_2328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5528_ (.X(_2329_),
    .A(_2310_),
    .B(_2313_),
    .C(_2328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5529_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2310_),
    .A2(_2313_),
    .Y(_2330_),
    .B1(_2328_));
 sg13g2_o21ai_1 _5530_ (.B1(net592),
    .VDD(VPWR),
    .Y(_2331_),
    .VSS(VGND),
    .A1(_2329_),
    .A2(_2330_));
 sg13g2_o21ai_1 _5531_ (.B1(_2331_),
    .VDD(VPWR),
    .Y(_2332_),
    .VSS(VGND),
    .A1(net592),
    .A2(net1089));
 sg13g2_nor2_1 _5532_ (.A(net463),
    .B(_2332_),
    .Y(_0317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5533_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net520),
    .A2(\mydesign.pe_weights[23] ),
    .Y(_2333_),
    .B1(\mydesign.accum[14] ));
 sg13g2_nand3_1 _5534_ (.B(net520),
    .C(\mydesign.pe_weights[23] ),
    .A(\mydesign.accum[14] ),
    .Y(_2334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5535_ (.Y(_2335_),
    .B(_2334_),
    .A_N(_2333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5536_ (.B1(_2318_),
    .VDD(VPWR),
    .Y(_2336_),
    .VSS(VGND),
    .A1(_2316_),
    .A2(_2319_));
 sg13g2_inv_1 _5537_ (.VDD(VPWR),
    .Y(_2337_),
    .A(_2336_),
    .VSS(VGND));
 sg13g2_xnor2_1 _5538_ (.Y(_2338_),
    .A(_2335_),
    .B(_2336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5539_ (.B(_2322_),
    .C(_2338_),
    .A(_2321_),
    .Y(_2339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5540_ (.A2(_2322_),
    .A1(_2321_),
    .B1(_2338_),
    .X(_2340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5541_ (.A(_2339_),
    .B(_2340_),
    .X(_2341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5542_ (.B(_2324_),
    .C(_2341_),
    .A(_2323_),
    .Y(_2342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5543_ (.Y(_2343_),
    .A(_2325_),
    .B(_2341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5544_ (.A(_2327_),
    .B(_2330_),
    .C(_2343_),
    .Y(_2344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5545_ (.B1(_2343_),
    .VDD(VPWR),
    .Y(_2345_),
    .VSS(VGND),
    .A1(_2327_),
    .A2(_2330_));
 sg13g2_nand2b_1 _5546_ (.Y(_2346_),
    .B(_2345_),
    .A_N(_2344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5547_ (.B1(net481),
    .VDD(VPWR),
    .Y(_2347_),
    .VSS(VGND),
    .A1(net592),
    .A2(net1052));
 sg13g2_a21oi_1 _5548_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net592),
    .A2(_2346_),
    .Y(_0318_),
    .B1(_2347_));
 sg13g2_nand2_1 _5549_ (.Y(_2348_),
    .A(_2342_),
    .B(_2345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5550_ (.B1(_2334_),
    .VDD(VPWR),
    .Y(_2349_),
    .VSS(VGND),
    .A1(_2333_),
    .A2(_2337_));
 sg13g2_xnor2_1 _5551_ (.Y(_2350_),
    .A(\mydesign.accum[15] ),
    .B(_2349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5552_ (.Y(_2351_),
    .A(_2339_),
    .B(_2350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5553_ (.B(_2351_),
    .A(_2348_),
    .X(_2352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5554_ (.B1(net481),
    .VDD(VPWR),
    .Y(_2353_),
    .VSS(VGND),
    .A1(net592),
    .A2(net1055));
 sg13g2_a21oi_1 _5555_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net592),
    .A2(_2352_),
    .Y(_0319_),
    .B1(_2353_));
 sg13g2_nor2_2 _5556_ (.A(_2607_),
    .B(_2683_),
    .Y(_2354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _5557_ (.Y(_2355_),
    .A(net606),
    .B(_2354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _5558_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net608),
    .Y(_2356_),
    .A2(_2354_),
    .A1(net606));
 sg13g2_nand2_1 _5559_ (.Y(_2357_),
    .A(net416),
    .B(_2356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5560_ (.B1(_2357_),
    .VDD(VPWR),
    .Y(_0320_),
    .VSS(VGND),
    .A1(net603),
    .A2(_2355_));
 sg13g2_nand2_1 _5561_ (.Y(_2358_),
    .A(net658),
    .B(_2356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5562_ (.B1(_2358_),
    .VDD(VPWR),
    .Y(_0321_),
    .VSS(VGND),
    .A1(net601),
    .A2(_2355_));
 sg13g2_nand2_1 _5563_ (.Y(_2359_),
    .A(net650),
    .B(_2356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5564_ (.B1(_2359_),
    .VDD(VPWR),
    .Y(_0322_),
    .VSS(VGND),
    .A1(net599),
    .A2(_2355_));
 sg13g2_nand2_1 _5565_ (.Y(_2360_),
    .A(net680),
    .B(_2356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5566_ (.B1(_2360_),
    .VDD(VPWR),
    .Y(_0323_),
    .VSS(VGND),
    .A1(net597),
    .A2(_2355_));
 sg13g2_and3_1 _5567_ (.X(_2361_),
    .A(net587),
    .B(\mydesign.pe_inputs[4] ),
    .C(\mydesign.pe_weights[16] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5568_ (.B1(net475),
    .VDD(VPWR),
    .Y(_2362_),
    .VSS(VGND),
    .A1(net749),
    .A2(_2361_));
 sg13g2_a21oi_1 _5569_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net749),
    .A2(_2361_),
    .Y(_0324_),
    .B1(_2362_));
 sg13g2_nand2_1 _5570_ (.Y(_2363_),
    .A(\mydesign.pe_inputs[4] ),
    .B(\mydesign.pe_weights[17] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5571_ (.X(_2364_),
    .A(\mydesign.accum[1] ),
    .B(\mydesign.pe_inputs[5] ),
    .C(net523),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5572_ (.B(\mydesign.pe_inputs[5] ),
    .C(net524),
    .A(\mydesign.accum[1] ),
    .Y(_2365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5573_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_inputs[5] ),
    .A2(net524),
    .Y(_2366_),
    .B1(\mydesign.accum[1] ));
 sg13g2_nor2_1 _5574_ (.A(_2364_),
    .B(_2366_),
    .Y(_2367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5575_ (.Y(_2368_),
    .A(_2363_),
    .B(_2367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5576_ (.B(\mydesign.pe_inputs[4] ),
    .C(net524),
    .A(net749),
    .Y(_2369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5577_ (.A(net749),
    .B(\mydesign.pe_inputs[4] ),
    .C(net523),
    .D(_2368_),
    .X(_2370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5578_ (.B(_2369_),
    .A(_2368_),
    .X(_2371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5579_ (.B1(net475),
    .VDD(VPWR),
    .Y(_2372_),
    .VSS(VGND),
    .A1(net587),
    .A2(net1057));
 sg13g2_a21oi_1 _5580_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net587),
    .A2(_2371_),
    .Y(_0325_),
    .B1(_2372_));
 sg13g2_nand2_1 _5581_ (.Y(_2373_),
    .A(\mydesign.pe_inputs[4] ),
    .B(net1017),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5582_ (.B1(_2365_),
    .VDD(VPWR),
    .Y(_2374_),
    .VSS(VGND),
    .A1(_2363_),
    .A2(_2366_));
 sg13g2_nand2_1 _5583_ (.Y(_2375_),
    .A(\mydesign.pe_inputs[5] ),
    .B(\mydesign.pe_weights[17] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5584_ (.X(_2376_),
    .A(\mydesign.accum[2] ),
    .B(\mydesign.pe_inputs[6] ),
    .C(net523),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5585_ (.B(\mydesign.pe_inputs[6] ),
    .C(net523),
    .A(\mydesign.accum[2] ),
    .Y(_2377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5586_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.pe_inputs[6] ),
    .A2(net523),
    .Y(_2378_),
    .B1(\mydesign.accum[2] ));
 sg13g2_nor2_1 _5587_ (.A(_2376_),
    .B(_2378_),
    .Y(_2379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5588_ (.Y(_2380_),
    .A(_2375_),
    .B(_2379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5589_ (.Y(_2381_),
    .A(_2374_),
    .B(_2380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5590_ (.Y(_2382_),
    .A(_2374_),
    .B(_2380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5591_ (.B(_2382_),
    .A(_2373_),
    .X(_2383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5592_ (.Y(_2384_),
    .A(_2370_),
    .B(_2383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5593_ (.Y(_2385_),
    .A(_2370_),
    .B(_2383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5594_ (.B1(net476),
    .VDD(VPWR),
    .Y(_2386_),
    .VSS(VGND),
    .A1(net586),
    .A2(net1040));
 sg13g2_a21oi_1 _5595_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net586),
    .A2(_2385_),
    .Y(_0326_),
    .B1(_2386_));
 sg13g2_nand2_1 _5596_ (.Y(_2387_),
    .A(net1111),
    .B(\mydesign.pe_weights[19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5597_ (.B1(_2381_),
    .VDD(VPWR),
    .Y(_2388_),
    .VSS(VGND),
    .A1(_2373_),
    .A2(_2382_));
 sg13g2_nand2_1 _5598_ (.Y(_2389_),
    .A(\mydesign.pe_inputs[5] ),
    .B(\mydesign.pe_weights[18] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5599_ (.B1(_2377_),
    .VDD(VPWR),
    .Y(_2390_),
    .VSS(VGND),
    .A1(_2375_),
    .A2(_2378_));
 sg13g2_nand2_1 _5600_ (.Y(_2391_),
    .A(\mydesign.pe_inputs[6] ),
    .B(\mydesign.pe_weights[17] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5601_ (.X(_2392_),
    .A(\mydesign.accum[3] ),
    .B(net519),
    .C(net523),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5602_ (.B(\mydesign.pe_inputs[7] ),
    .C(net523),
    .A(\mydesign.accum[3] ),
    .Y(_2393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5603_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net519),
    .A2(net523),
    .Y(_2394_),
    .B1(\mydesign.accum[3] ));
 sg13g2_nor2_1 _5604_ (.A(_2392_),
    .B(_2394_),
    .Y(_2395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5605_ (.Y(_2396_),
    .A(_2391_),
    .B(_2395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5606_ (.Y(_2397_),
    .A(_2390_),
    .B(_2396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5607_ (.A(_2390_),
    .B(_2396_),
    .Y(_2398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5608_ (.B(_2396_),
    .A(_2390_),
    .X(_2399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5609_ (.Y(_2400_),
    .A(_2389_),
    .B(_2399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5610_ (.Y(_2401_),
    .A(_2388_),
    .B(_2400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5611_ (.Y(_2402_),
    .A(_2388_),
    .B(_2400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5612_ (.B(_2402_),
    .A(_2387_),
    .X(_2403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5613_ (.Y(_2404_),
    .B(_2403_),
    .A_N(_2384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5614_ (.B(_2403_),
    .A(_2384_),
    .X(_2405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5615_ (.B1(net476),
    .VDD(VPWR),
    .Y(_2406_),
    .VSS(VGND),
    .A1(net586),
    .A2(net1045));
 sg13g2_a21oi_1 _5616_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net586),
    .A2(_2405_),
    .Y(_0327_),
    .B1(_2406_));
 sg13g2_o21ai_1 _5617_ (.B1(_2401_),
    .VDD(VPWR),
    .Y(_2407_),
    .VSS(VGND),
    .A1(_2387_),
    .A2(_2402_));
 sg13g2_nand2_1 _5618_ (.Y(_2408_),
    .A(\mydesign.pe_inputs[5] ),
    .B(\mydesign.pe_weights[19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5619_ (.B1(_2397_),
    .VDD(VPWR),
    .Y(_2409_),
    .VSS(VGND),
    .A1(_2389_),
    .A2(_2398_));
 sg13g2_nand2_1 _5620_ (.Y(_2410_),
    .A(\mydesign.pe_inputs[6] ),
    .B(\mydesign.pe_weights[18] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5621_ (.B(net519),
    .C(\mydesign.pe_weights[17] ),
    .A(\mydesign.accum[4] ),
    .Y(_2411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5622_ (.A2(\mydesign.pe_weights[17] ),
    .A1(net519),
    .B1(\mydesign.accum[4] ),
    .X(_2412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5623_ (.Y(_2413_),
    .A(_2411_),
    .B(_2412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5624_ (.B1(_2393_),
    .VDD(VPWR),
    .Y(_2414_),
    .VSS(VGND),
    .A1(_2391_),
    .A2(_2394_));
 sg13g2_inv_1 _5625_ (.VDD(VPWR),
    .Y(_2415_),
    .A(_2414_),
    .VSS(VGND));
 sg13g2_xnor2_1 _5626_ (.Y(_2416_),
    .A(_2413_),
    .B(_2414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5627_ (.Y(_2417_),
    .B(_2416_),
    .A_N(_2410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5628_ (.Y(_2418_),
    .A(_2410_),
    .B(_2416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5629_ (.Y(_2419_),
    .A(_2409_),
    .B(_2418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5630_ (.A(_2409_),
    .B(_2418_),
    .Y(_2420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5631_ (.B(_2418_),
    .A(_2409_),
    .X(_2421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5632_ (.Y(_2422_),
    .A(_2408_),
    .B(_2421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5633_ (.Y(_2423_),
    .A(_2407_),
    .B(_2422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5634_ (.Y(_2424_),
    .A(_2407_),
    .B(_2422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5635_ (.Y(_2425_),
    .A(_2404_),
    .B(_2424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5636_ (.B1(net476),
    .VDD(VPWR),
    .Y(_2426_),
    .VSS(VGND),
    .A1(net586),
    .A2(net1068));
 sg13g2_a21oi_1 _5637_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net586),
    .A2(_2425_),
    .Y(_0328_),
    .B1(_2426_));
 sg13g2_o21ai_1 _5638_ (.B1(_2423_),
    .VDD(VPWR),
    .Y(_2427_),
    .VSS(VGND),
    .A1(_2404_),
    .A2(_2424_));
 sg13g2_o21ai_1 _5639_ (.B1(_2419_),
    .VDD(VPWR),
    .Y(_2428_),
    .VSS(VGND),
    .A1(_2408_),
    .A2(_2420_));
 sg13g2_nand2_1 _5640_ (.Y(_2429_),
    .A(\mydesign.pe_inputs[6] ),
    .B(\mydesign.pe_weights[19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5641_ (.B1(_2417_),
    .VDD(VPWR),
    .Y(_2430_),
    .VSS(VGND),
    .A1(_2413_),
    .A2(_2415_));
 sg13g2_nand4_1 _5642_ (.B(\mydesign.accum[4] ),
    .C(net519),
    .A(\mydesign.accum[5] ),
    .Y(_2431_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\mydesign.pe_weights[17] ));
 sg13g2_xor2_1 _5643_ (.B(_2411_),
    .A(\mydesign.accum[5] ),
    .X(_2432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5644_ (.Y(_2433_),
    .A(net519),
    .B(\mydesign.pe_weights[18] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5645_ (.B(_2433_),
    .A(_2432_),
    .X(_2434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5646_ (.Y(_2435_),
    .A(_2430_),
    .B(_2434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5647_ (.A(_2430_),
    .B(_2434_),
    .Y(_2436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5648_ (.B(_2434_),
    .A(_2430_),
    .X(_2437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5649_ (.Y(_2438_),
    .A(_2429_),
    .B(_2437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5650_ (.Y(_2439_),
    .A(_2428_),
    .B(_2438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5651_ (.B(_2438_),
    .A(_2428_),
    .X(_2440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5652_ (.Y(_2441_),
    .A(_2427_),
    .B(_2440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5653_ (.Y(_2442_),
    .A(_2427_),
    .B(_2440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5654_ (.B1(net476),
    .VDD(VPWR),
    .Y(_2443_),
    .VSS(VGND),
    .A1(net586),
    .A2(net1063));
 sg13g2_a21oi_1 _5655_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net586),
    .A2(_2442_),
    .Y(_0329_),
    .B1(_2443_));
 sg13g2_o21ai_1 _5656_ (.B1(_2435_),
    .VDD(VPWR),
    .Y(_2444_),
    .VSS(VGND),
    .A1(_2429_),
    .A2(_2436_));
 sg13g2_o21ai_1 _5657_ (.B1(_2431_),
    .VDD(VPWR),
    .Y(_2445_),
    .VSS(VGND),
    .A1(_2432_),
    .A2(_2433_));
 sg13g2_xor2_1 _5658_ (.B(_2445_),
    .A(\mydesign.accum[6] ),
    .X(_2446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5659_ (.X(_2447_),
    .A(net519),
    .B(\mydesign.pe_weights[19] ),
    .C(_2446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5660_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net519),
    .A2(\mydesign.pe_weights[19] ),
    .Y(_2448_),
    .B1(_2446_));
 sg13g2_or2_1 _5661_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2449_),
    .B(_2448_),
    .A(_2447_));
 sg13g2_inv_1 _5662_ (.VDD(VPWR),
    .Y(_2450_),
    .A(_2449_),
    .VSS(VGND));
 sg13g2_xnor2_1 _5663_ (.Y(_2451_),
    .A(_2444_),
    .B(_2450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5664_ (.X(_2452_),
    .A(_2439_),
    .B(_2441_),
    .C(_2451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5665_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2439_),
    .A2(_2441_),
    .Y(_2453_),
    .B1(_2451_));
 sg13g2_or2_1 _5666_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2454_),
    .B(_2453_),
    .A(_2452_));
 sg13g2_o21ai_1 _5667_ (.B1(net476),
    .VDD(VPWR),
    .Y(_2455_),
    .VSS(VGND),
    .A1(net587),
    .A2(net1049));
 sg13g2_a21oi_1 _5668_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net587),
    .A2(_2454_),
    .Y(_0330_),
    .B1(_2455_));
 sg13g2_a21oi_1 _5669_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mydesign.accum[6] ),
    .A2(_2445_),
    .Y(_2456_),
    .B1(_2447_));
 sg13g2_a21oi_1 _5670_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2444_),
    .A2(_2450_),
    .Y(_2457_),
    .B1(_2453_));
 sg13g2_o21ai_1 _5671_ (.B1(net587),
    .VDD(VPWR),
    .Y(_2458_),
    .VSS(VGND),
    .A1(_2456_),
    .A2(_2457_));
 sg13g2_a21oi_2 _5672_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2458_),
    .Y(_2459_),
    .A2(_2457_),
    .A1(_2456_));
 sg13g2_o21ai_1 _5673_ (.B1(net473),
    .VDD(VPWR),
    .Y(_2460_),
    .VSS(VGND),
    .A1(net409),
    .A2(_2459_));
 sg13g2_a21oi_1 _5674_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net409),
    .A2(_2459_),
    .Y(_0331_),
    .B1(_2460_));
 sg13g2_nand2_2 _5675_ (.Y(_2461_),
    .A(net462),
    .B(_2684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5676_ (.Y(_2462_),
    .A(net683),
    .B(_2461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5677_ (.B1(_2462_),
    .VDD(VPWR),
    .Y(_0332_),
    .VSS(VGND),
    .A1(net604),
    .A2(_2461_));
 sg13g2_nand2_1 _5678_ (.Y(_2463_),
    .A(net679),
    .B(_2461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5679_ (.B1(_2463_),
    .VDD(VPWR),
    .Y(_0333_),
    .VSS(VGND),
    .A1(net602),
    .A2(_2461_));
 sg13g2_nand2_1 _5680_ (.Y(_2464_),
    .A(net645),
    .B(_2461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5681_ (.B1(_2464_),
    .VDD(VPWR),
    .Y(_0334_),
    .VSS(VGND),
    .A1(net600),
    .A2(_2461_));
 sg13g2_nand2_1 _5682_ (.Y(_2465_),
    .A(net649),
    .B(_2461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5683_ (.B1(_2465_),
    .VDD(VPWR),
    .Y(_0335_),
    .VSS(VGND),
    .A1(net598),
    .A2(_2461_));
 sg13g2_nand3_1 _5684_ (.B(_2599_),
    .C(_0384_),
    .A(net618),
    .Y(_2466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5685_ (.A(net608),
    .B(_2698_),
    .Y(_2467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5686_ (.Y(_2468_),
    .A(net623),
    .B(net430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5687_ (.Y(_2469_),
    .A(net755),
    .B(_2466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5688_ (.B1(_2469_),
    .VDD(VPWR),
    .Y(_0336_),
    .VSS(VGND),
    .A1(net755),
    .A2(_2468_));
 sg13g2_nor3_1 _5689_ (.A(net457),
    .B(net456),
    .C(_2468_),
    .Y(_2470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5690_ (.A2(_2466_),
    .A1(net834),
    .B1(_2470_),
    .X(_0337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5691_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net512),
    .A2(net457),
    .Y(_2471_),
    .B1(_2468_));
 sg13g2_nor2_1 _5692_ (.A(_2466_),
    .B(_2471_),
    .Y(_2472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5693_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net457),
    .A2(_2467_),
    .Y(_2473_),
    .B1(net512));
 sg13g2_nor2_1 _5694_ (.A(_2472_),
    .B(_2473_),
    .Y(_0338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5695_ (.B(net457),
    .C(_2467_),
    .A(net512),
    .Y(_2474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5696_ (.B1(net504),
    .VDD(VPWR),
    .Y(_2475_),
    .VSS(VGND),
    .A1(_2466_),
    .A2(_2471_));
 sg13g2_o21ai_1 _5697_ (.B1(_2475_),
    .VDD(VPWR),
    .Y(_0339_),
    .VSS(VGND),
    .A1(net504),
    .A2(_2474_));
 sg13g2_nand3_1 _5698_ (.B(net610),
    .C(_2656_),
    .A(\mydesign.load_counter[3] ),
    .Y(_2476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5699_ (.B(net725),
    .C(_2476_),
    .A(net613),
    .Y(_2477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5700_ (.B1(_2477_),
    .VDD(VPWR),
    .Y(_0340_),
    .VSS(VGND),
    .A1(net603),
    .A2(_2476_));
 sg13g2_nand3_1 _5701_ (.B(net717),
    .C(_2476_),
    .A(net613),
    .Y(_2478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5702_ (.B1(_2478_),
    .VDD(VPWR),
    .Y(_0341_),
    .VSS(VGND),
    .A1(net601),
    .A2(_2476_));
 sg13g2_nand3_1 _5703_ (.B(net705),
    .C(_2476_),
    .A(net613),
    .Y(_2479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5704_ (.B1(_2479_),
    .VDD(VPWR),
    .Y(_0342_),
    .VSS(VGND),
    .A1(net599),
    .A2(_2476_));
 sg13g2_nand3_1 _5705_ (.B(net731),
    .C(_2476_),
    .A(net613),
    .Y(_2480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5706_ (.B1(_2480_),
    .VDD(VPWR),
    .Y(_0343_),
    .VSS(VGND),
    .A1(net597),
    .A2(_2476_));
 sg13g2_a21o_2 _5707_ (.A2(_2354_),
    .A1(net610),
    .B1(net609),
    .X(_2481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5708_ (.A(_2605_),
    .B(_2639_),
    .C(_2683_),
    .Y(_2482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5709_ (.A(\mydesign.load_counter[1] ),
    .B(_2605_),
    .C(_2607_),
    .Y(_2483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _5710_ (.A(net432),
    .B(_2482_),
    .C(_2483_),
    .Y(_2484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _5711_ (.A(_2520_),
    .B(_2484_),
    .Y(_2485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5712_ (.A0(net802),
    .A1(_2485_),
    .S(_2481_),
    .X(_0344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _5713_ (.A(_2519_),
    .B(_2484_),
    .Y(_2486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5714_ (.A0(net774),
    .A1(_2486_),
    .S(_2481_),
    .X(_0345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _5715_ (.A(_2518_),
    .B(_2484_),
    .Y(_2487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5716_ (.A0(net770),
    .A1(_2487_),
    .S(_2481_),
    .X(_0346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _5717_ (.A(_2517_),
    .B(_2484_),
    .Y(_2488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5718_ (.A0(net777),
    .A1(_2488_),
    .S(_2481_),
    .X(_0347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _5719_ (.Y(_2489_),
    .B(net614),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2482_));
 sg13g2_mux2_1 _5720_ (.A0(net771),
    .A1(_2485_),
    .S(_2489_),
    .X(_0348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5721_ (.A0(net764),
    .A1(_2486_),
    .S(_2489_),
    .X(_0349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5722_ (.A0(net761),
    .A1(_2487_),
    .S(_2489_),
    .X(_0350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5723_ (.A0(net763),
    .A1(_2488_),
    .S(_2489_),
    .X(_0351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5724_ (.B(_2619_),
    .C(_2621_),
    .A(net611),
    .Y(_2490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5725_ (.B(net723),
    .C(_2490_),
    .A(net615),
    .Y(_2491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5726_ (.B1(_2491_),
    .VDD(VPWR),
    .Y(_0352_),
    .VSS(VGND),
    .A1(net604),
    .A2(_2490_));
 sg13g2_nand3_1 _5727_ (.B(net716),
    .C(_2490_),
    .A(net615),
    .Y(_2492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5728_ (.B1(_2492_),
    .VDD(VPWR),
    .Y(_0353_),
    .VSS(VGND),
    .A1(net602),
    .A2(_2490_));
 sg13g2_nand3_1 _5729_ (.B(net711),
    .C(_2490_),
    .A(net615),
    .Y(_2493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5730_ (.B1(_2493_),
    .VDD(VPWR),
    .Y(_0354_),
    .VSS(VGND),
    .A1(net600),
    .A2(_2490_));
 sg13g2_nand3_1 _5731_ (.B(net714),
    .C(_2490_),
    .A(net620),
    .Y(_2494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5732_ (.B1(_2494_),
    .VDD(VPWR),
    .Y(_0355_),
    .VSS(VGND),
    .A1(net598),
    .A2(_2490_));
 sg13g2_nand2_2 _5733_ (.Y(_2495_),
    .A(net462),
    .B(_2686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5734_ (.Y(_2496_),
    .A(net647),
    .B(_2495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5735_ (.B1(_2496_),
    .VDD(VPWR),
    .Y(_0356_),
    .VSS(VGND),
    .A1(net604),
    .A2(_2495_));
 sg13g2_nand2_1 _5736_ (.Y(_2497_),
    .A(net700),
    .B(_2495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5737_ (.B1(_2497_),
    .VDD(VPWR),
    .Y(_0357_),
    .VSS(VGND),
    .A1(net602),
    .A2(_2495_));
 sg13g2_nand2_1 _5738_ (.Y(_2498_),
    .A(net694),
    .B(_2495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5739_ (.B1(_2498_),
    .VDD(VPWR),
    .Y(_0358_),
    .VSS(VGND),
    .A1(net600),
    .A2(_2495_));
 sg13g2_nand2_1 _5740_ (.Y(_2499_),
    .A(net722),
    .B(_2495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5741_ (.B1(_2499_),
    .VDD(VPWR),
    .Y(_0359_),
    .VSS(VGND),
    .A1(net598),
    .A2(_2495_));
 sg13g2_o21ai_1 _5742_ (.B1(net462),
    .VDD(VPWR),
    .Y(_2500_),
    .VSS(VGND),
    .A1(net608),
    .A2(_2663_));
 sg13g2_nand2_1 _5743_ (.Y(_2501_),
    .A(net748),
    .B(_2500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5744_ (.B1(_2501_),
    .VDD(VPWR),
    .Y(_0360_),
    .VSS(VGND),
    .A1(_1769_),
    .A2(_2500_));
 sg13g2_nand2_1 _5745_ (.Y(_2502_),
    .A(net727),
    .B(_2500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5746_ (.B1(_2502_),
    .VDD(VPWR),
    .Y(_0361_),
    .VSS(VGND),
    .A1(_1771_),
    .A2(_2500_));
 sg13g2_nand2_1 _5747_ (.Y(_2503_),
    .A(net698),
    .B(_2500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5748_ (.B1(_2503_),
    .VDD(VPWR),
    .Y(_0362_),
    .VSS(VGND),
    .A1(_1773_),
    .A2(_2500_));
 sg13g2_nand2_1 _5749_ (.Y(_2504_),
    .A(net751),
    .B(_2500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5750_ (.B1(_2504_),
    .VDD(VPWR),
    .Y(_0363_),
    .VSS(VGND),
    .A1(_1775_),
    .A2(_2500_));
 sg13g2_nor3_2 _5751_ (.A(_2591_),
    .B(_2622_),
    .C(_2648_),
    .Y(_2505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5752_ (.B1(net612),
    .VDD(VPWR),
    .Y(_2506_),
    .VSS(VGND),
    .A1(net985),
    .A2(_2505_));
 sg13g2_a21oi_1 _5753_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1769_),
    .A2(_2505_),
    .Y(_0364_),
    .B1(net986));
 sg13g2_o21ai_1 _5754_ (.B1(net612),
    .VDD(VPWR),
    .Y(_2507_),
    .VSS(VGND),
    .A1(net823),
    .A2(_2505_));
 sg13g2_a21oi_1 _5755_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1771_),
    .A2(_2505_),
    .Y(_0365_),
    .B1(net824));
 sg13g2_o21ai_1 _5756_ (.B1(net612),
    .VDD(VPWR),
    .Y(_2508_),
    .VSS(VGND),
    .A1(net930),
    .A2(_2505_));
 sg13g2_a21oi_1 _5757_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1773_),
    .A2(_2505_),
    .Y(_0366_),
    .B1(net931));
 sg13g2_o21ai_1 _5758_ (.B1(net612),
    .VDD(VPWR),
    .Y(_2509_),
    .VSS(VGND),
    .A1(net869),
    .A2(_2505_));
 sg13g2_a21oi_1 _5759_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1775_),
    .A2(_2505_),
    .Y(_0367_),
    .B1(net870));
 sg13g2_o21ai_1 _5760_ (.B1(net615),
    .VDD(VPWR),
    .Y(_2510_),
    .VSS(VGND),
    .A1(_2591_),
    .A2(_1400_));
 sg13g2_mux2_1 _5761_ (.A0(net767),
    .A1(_2485_),
    .S(_2510_),
    .X(_0368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5762_ (.A0(net803),
    .A1(_2486_),
    .S(_2510_),
    .X(_0369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5763_ (.A0(net784),
    .A1(_2487_),
    .S(_2510_),
    .X(_0370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5764_ (.A0(net781),
    .A1(_2488_),
    .S(_2510_),
    .X(_0371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _5765_ (.Y(_2511_),
    .A(net462),
    .B(_0910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5766_ (.Y(_2512_),
    .A(net699),
    .B(_2511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5767_ (.B1(_2512_),
    .VDD(VPWR),
    .Y(_0372_),
    .VSS(VGND),
    .A1(net604),
    .A2(_2511_));
 sg13g2_nand2_1 _5768_ (.Y(_2513_),
    .A(net693),
    .B(_2511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5769_ (.B1(_2513_),
    .VDD(VPWR),
    .Y(_0373_),
    .VSS(VGND),
    .A1(net602),
    .A2(_2511_));
 sg13g2_nand2_1 _5770_ (.Y(_2514_),
    .A(net737),
    .B(_2511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5771_ (.B1(_2514_),
    .VDD(VPWR),
    .Y(_0374_),
    .VSS(VGND),
    .A1(net600),
    .A2(_2511_));
 sg13g2_nand2_1 _5772_ (.Y(_2515_),
    .A(net674),
    .B(_2511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5773_ (.B1(_2515_),
    .VDD(VPWR),
    .Y(_0375_),
    .VSS(VGND),
    .A1(net598),
    .A2(_2511_));
 sg13g2_dfrbpq_1 _5774_ (.RESET_B(net240),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0000_),
    .Q(\mydesign.valid_out ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _5775_ (.RESET_B(net183),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0001_),
    .Q(\mydesign.weights[2][4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5776_ (.RESET_B(net181),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0002_),
    .Q(\mydesign.weights[2][5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5777_ (.RESET_B(net179),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0003_),
    .Q(\mydesign.weights[2][6] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5778_ (.RESET_B(net177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net753),
    .Q(\mydesign.weights[2][7] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5779_ (.RESET_B(net175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0005_),
    .Q(\mydesign.inputs[0][24] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _5780_ (.RESET_B(net174),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0006_),
    .Q(\mydesign.inputs[0][25] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _5781_ (.RESET_B(net173),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0007_),
    .Q(\mydesign.inputs[0][26] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _5782_ (.RESET_B(net172),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0008_),
    .Q(\mydesign.inputs[0][27] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _5783_ (.RESET_B(net171),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net678),
    .Q(\mydesign.weights[2][16] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5784_ (.RESET_B(net169),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net676),
    .Q(\mydesign.weights[2][17] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5785_ (.RESET_B(net167),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0011_),
    .Q(\mydesign.weights[2][18] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5786_ (.RESET_B(net165),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net663),
    .Q(\mydesign.weights[2][19] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5787_ (.RESET_B(net163),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net424),
    .Q(\mydesign.inputs[2][8] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _5788_ (.RESET_B(net162),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net421),
    .Q(\mydesign.inputs[2][9] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5789_ (.RESET_B(net161),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net668),
    .Q(\mydesign.inputs[2][10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _5790_ (.RESET_B(net160),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net643),
    .Q(\mydesign.inputs[2][11] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5791_ (.RESET_B(net159),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0017_),
    .Q(\mydesign.inputs[2][4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _5792_ (.RESET_B(net158),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0018_),
    .Q(\mydesign.inputs[2][5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _5793_ (.RESET_B(net157),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0019_),
    .Q(\mydesign.inputs[2][6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _5794_ (.RESET_B(net156),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0020_),
    .Q(\mydesign.inputs[2][7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _5795_ (.RESET_B(net155),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0021_),
    .Q(\mydesign.inputs[1][8] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _5796_ (.RESET_B(net154),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0022_),
    .Q(\mydesign.inputs[1][9] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _5797_ (.RESET_B(net153),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0023_),
    .Q(\mydesign.inputs[1][10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _5798_ (.RESET_B(net152),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0024_),
    .Q(\mydesign.inputs[1][11] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _5799_ (.RESET_B(net151),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0025_),
    .Q(\mydesign.inputs[1][12] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _5800_ (.RESET_B(net150),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0026_),
    .Q(\mydesign.inputs[1][13] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5801_ (.RESET_B(net149),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0027_),
    .Q(\mydesign.inputs[1][14] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5802_ (.RESET_B(net148),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0028_),
    .Q(\mydesign.inputs[1][15] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5803_ (.RESET_B(net147),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0029_),
    .Q(\mydesign.weights[2][12] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5804_ (.RESET_B(net145),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0030_),
    .Q(\mydesign.weights[2][13] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5805_ (.RESET_B(net143),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0031_),
    .Q(\mydesign.weights[2][14] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5806_ (.RESET_B(net141),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0032_),
    .Q(\mydesign.weights[2][15] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5807_ (.RESET_B(net139),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0033_),
    .Q(\mydesign.inputs[2][16] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5808_ (.RESET_B(net137),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0034_),
    .Q(\mydesign.inputs[2][17] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5809_ (.RESET_B(net135),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0035_),
    .Q(\mydesign.inputs[2][18] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5810_ (.RESET_B(net133),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0036_),
    .Q(\mydesign.inputs[2][19] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5811_ (.RESET_B(net131),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0037_),
    .Q(\mydesign.inputs[1][16] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _5812_ (.RESET_B(net130),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0038_),
    .Q(\mydesign.inputs[1][17] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5813_ (.RESET_B(net129),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0039_),
    .Q(\mydesign.inputs[1][18] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5814_ (.RESET_B(net128),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0040_),
    .Q(\mydesign.inputs[1][19] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _5815_ (.RESET_B(net127),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0041_),
    .Q(\mydesign.inputs[1][20] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _5816_ (.RESET_B(net126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0042_),
    .Q(\mydesign.inputs[1][21] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5817_ (.RESET_B(net125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0043_),
    .Q(\mydesign.inputs[1][22] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5818_ (.RESET_B(net124),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0044_),
    .Q(\mydesign.inputs[1][23] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _5819_ (.RESET_B(net123),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0045_),
    .Q(\mydesign.inputs[0][12] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _5820_ (.RESET_B(net122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0046_),
    .Q(\mydesign.inputs[0][13] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5821_ (.RESET_B(net121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0047_),
    .Q(\mydesign.inputs[0][14] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5822_ (.RESET_B(net120),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0048_),
    .Q(\mydesign.inputs[0][15] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5823_ (.RESET_B(net119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0049_),
    .Q(\mydesign.inputs[0][16] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _5824_ (.RESET_B(net118),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0050_),
    .Q(\mydesign.inputs[0][17] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5825_ (.RESET_B(net117),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0051_),
    .Q(\mydesign.inputs[0][18] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5826_ (.RESET_B(net116),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0052_),
    .Q(\mydesign.inputs[0][19] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5827_ (.RESET_B(net115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net710),
    .Q(\mydesign.inputs[3][0] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _5828_ (.RESET_B(net113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net743),
    .Q(\mydesign.inputs[3][1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _5829_ (.RESET_B(net111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net713),
    .Q(\mydesign.inputs[3][2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _5830_ (.RESET_B(net109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net720),
    .Q(\mydesign.inputs[3][3] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _5831_ (.RESET_B(net107),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0057_),
    .Q(\mydesign.load_counter[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5832_ (.RESET_B(net105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0058_),
    .Q(\mydesign.load_counter[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5833_ (.RESET_B(net103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0059_),
    .Q(\mydesign.load_counter[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5834_ (.RESET_B(net101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0060_),
    .Q(\mydesign.load_counter[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5835_ (.RESET_B(net99),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0061_),
    .Q(\mydesign.compute_en ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _5836_ (.RESET_B(net97),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0062_),
    .Q(\mydesign.cp[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5837_ (.RESET_B(net95),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0063_),
    .Q(\mydesign.cp[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5838_ (.RESET_B(net93),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0064_),
    .Q(\mydesign.cp[2] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _5839_ (.RESET_B(net91),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0065_),
    .Q(\mydesign.cp2[0] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _5840_ (.RESET_B(net89),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0066_),
    .Q(\mydesign.cp2[1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _5841_ (.RESET_B(net87),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net408),
    .Q(\mydesign.cp2[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _5842_ (.RESET_B(net85),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0068_),
    .Q(net8),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5843_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1070),
    .Q(net9),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _5844_ (.RESET_B(net81),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0070_),
    .Q(net10),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _5845_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0071_),
    .Q(net11),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _5846_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0072_),
    .Q(net12),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _5847_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0073_),
    .Q(net13),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _5848_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0074_),
    .Q(net14),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5849_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1085),
    .Q(net15),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5850_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net415),
    .Q(\mydesign.inputs[2][12] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5851_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net426),
    .Q(\mydesign.inputs[2][13] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5852_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net419),
    .Q(\mydesign.inputs[2][14] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5853_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net653),
    .Q(\mydesign.inputs[2][15] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _5854_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0080_),
    .Q(\mydesign.pe_inputs[60] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _5855_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0081_),
    .Q(\mydesign.pe_inputs[61] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5856_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0082_),
    .Q(\mydesign.pe_inputs[62] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _5857_ (.RESET_B(net59),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0083_),
    .Q(\mydesign.pe_inputs[63] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5858_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net809),
    .Q(\mydesign.pe_weights[60] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5859_ (.RESET_B(net55),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0085_),
    .Q(\mydesign.pe_weights[61] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5860_ (.RESET_B(net53),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0086_),
    .Q(\mydesign.pe_weights[62] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5861_ (.RESET_B(net51),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0087_),
    .Q(\mydesign.pe_weights[63] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _5862_ (.RESET_B(net49),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0088_),
    .Q(\mydesign.accum[120] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5863_ (.RESET_B(net47),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0089_),
    .Q(\mydesign.accum[121] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5864_ (.RESET_B(net45),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0090_),
    .Q(\mydesign.accum[122] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5865_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0091_),
    .Q(\mydesign.accum[123] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5866_ (.RESET_B(net41),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0092_),
    .Q(\mydesign.accum[124] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5867_ (.RESET_B(net39),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0093_),
    .Q(\mydesign.accum[125] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5868_ (.RESET_B(net37),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0094_),
    .Q(\mydesign.accum[126] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5869_ (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0095_),
    .Q(\mydesign.accum[127] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5870_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1074),
    .Q(\mydesign.pe_inputs[56] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _5871_ (.RESET_B(net31),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1016),
    .Q(\mydesign.pe_inputs[57] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _5872_ (.RESET_B(net29),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1028),
    .Q(\mydesign.pe_inputs[58] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5873_ (.RESET_B(net27),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0099_),
    .Q(\mydesign.pe_inputs[59] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5874_ (.RESET_B(net25),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0100_),
    .Q(\mydesign.pe_weights[56] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5875_ (.RESET_B(net23),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0101_),
    .Q(\mydesign.pe_weights[57] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _5876_ (.RESET_B(net397),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0102_),
    .Q(\mydesign.pe_weights[58] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _5877_ (.RESET_B(net395),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0103_),
    .Q(\mydesign.pe_weights[59] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _5878_ (.RESET_B(net393),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0104_),
    .Q(\mydesign.accum[112] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _5879_ (.RESET_B(net391),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net852),
    .Q(\mydesign.accum[113] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _5880_ (.RESET_B(net389),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net878),
    .Q(\mydesign.accum[114] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5881_ (.RESET_B(net387),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0107_),
    .Q(\mydesign.accum[115] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5882_ (.RESET_B(net385),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0108_),
    .Q(\mydesign.accum[116] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5883_ (.RESET_B(net383),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0109_),
    .Q(\mydesign.accum[117] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _5884_ (.RESET_B(net381),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0110_),
    .Q(\mydesign.accum[118] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _5885_ (.RESET_B(net379),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0111_),
    .Q(\mydesign.accum[119] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5886_ (.RESET_B(net377),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net412),
    .Q(\mydesign.weights[3][4] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _5887_ (.RESET_B(net376),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net673),
    .Q(\mydesign.weights[3][5] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _5888_ (.RESET_B(net375),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net702),
    .Q(\mydesign.weights[3][6] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _5889_ (.RESET_B(net374),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net708),
    .Q(\mydesign.weights[3][7] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _5890_ (.RESET_B(net373),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0116_),
    .Q(\mydesign.pe_inputs[52] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _5891_ (.RESET_B(net371),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0117_),
    .Q(\mydesign.pe_inputs[53] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _5892_ (.RESET_B(net369),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0118_),
    .Q(\mydesign.pe_inputs[54] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _5893_ (.RESET_B(net367),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1047),
    .Q(\mydesign.pe_inputs[55] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _5894_ (.RESET_B(net365),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0120_),
    .Q(\mydesign.pe_weights[52] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _5895_ (.RESET_B(net363),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0121_),
    .Q(\mydesign.pe_weights[53] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _5896_ (.RESET_B(net361),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0122_),
    .Q(\mydesign.pe_weights[54] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _5897_ (.RESET_B(net359),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0123_),
    .Q(\mydesign.pe_weights[55] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _5898_ (.RESET_B(net357),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net689),
    .Q(\mydesign.accum[104] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _5899_ (.RESET_B(net355),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net917),
    .Q(\mydesign.accum[105] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _5900_ (.RESET_B(net353),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1011),
    .Q(\mydesign.accum[106] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _5901_ (.RESET_B(net351),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0127_),
    .Q(\mydesign.accum[107] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _5902_ (.RESET_B(net349),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0128_),
    .Q(\mydesign.accum[108] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _5903_ (.RESET_B(net347),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0129_),
    .Q(\mydesign.accum[109] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _5904_ (.RESET_B(net345),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0130_),
    .Q(\mydesign.accum[110] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _5905_ (.RESET_B(net343),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0131_),
    .Q(\mydesign.accum[111] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _5906_ (.RESET_B(net341),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0132_),
    .Q(\mydesign.inputs[0][20] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _5907_ (.RESET_B(net340),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0133_),
    .Q(\mydesign.inputs[0][21] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5908_ (.RESET_B(net339),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0134_),
    .Q(\mydesign.inputs[0][22] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5909_ (.RESET_B(net338),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0135_),
    .Q(\mydesign.inputs[0][23] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _5910_ (.RESET_B(net337),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0136_),
    .Q(\mydesign.pe_weights[48] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _5911_ (.RESET_B(net335),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0137_),
    .Q(\mydesign.pe_weights[49] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _5912_ (.RESET_B(net333),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0138_),
    .Q(\mydesign.pe_weights[50] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _5913_ (.RESET_B(net331),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0139_),
    .Q(\mydesign.pe_weights[51] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _5914_ (.RESET_B(net329),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0140_),
    .Q(\mydesign.accum[96] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _5915_ (.RESET_B(net327),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1008),
    .Q(\mydesign.accum[97] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _5916_ (.RESET_B(net325),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net848),
    .Q(\mydesign.accum[98] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _5917_ (.RESET_B(net323),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0143_),
    .Q(\mydesign.accum[99] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _5918_ (.RESET_B(net321),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0144_),
    .Q(\mydesign.accum[100] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _5919_ (.RESET_B(net319),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0145_),
    .Q(\mydesign.accum[101] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _5920_ (.RESET_B(net317),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0146_),
    .Q(\mydesign.accum[102] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _5921_ (.RESET_B(net315),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0147_),
    .Q(\mydesign.accum[103] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _5922_ (.RESET_B(net313),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0148_),
    .Q(\mydesign.pe_inputs[44] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5923_ (.RESET_B(net311),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0149_),
    .Q(\mydesign.pe_inputs[45] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5924_ (.RESET_B(net309),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0150_),
    .Q(\mydesign.pe_inputs[46] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5925_ (.RESET_B(net307),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0151_),
    .Q(\mydesign.pe_inputs[47] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5926_ (.RESET_B(net305),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0152_),
    .Q(\mydesign.pe_weights[44] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5927_ (.RESET_B(net303),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0153_),
    .Q(\mydesign.pe_weights[45] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5928_ (.RESET_B(net301),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net839),
    .Q(\mydesign.pe_weights[46] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _5929_ (.RESET_B(net299),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0155_),
    .Q(\mydesign.pe_weights[47] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _5930_ (.RESET_B(net297),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0156_),
    .Q(\mydesign.accum[88] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5931_ (.RESET_B(net295),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net897),
    .Q(\mydesign.accum[89] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _5932_ (.RESET_B(net293),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net965),
    .Q(\mydesign.accum[90] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _5933_ (.RESET_B(net291),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0159_),
    .Q(\mydesign.accum[91] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _5934_ (.RESET_B(net289),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0160_),
    .Q(\mydesign.accum[92] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _5935_ (.RESET_B(net287),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0161_),
    .Q(\mydesign.accum[93] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _5936_ (.RESET_B(net285),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0162_),
    .Q(\mydesign.accum[94] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5937_ (.RESET_B(net283),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0163_),
    .Q(\mydesign.accum[95] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5938_ (.RESET_B(net281),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1051),
    .Q(\mydesign.pe_inputs[40] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _5939_ (.RESET_B(net279),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0165_),
    .Q(\mydesign.pe_inputs[41] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _5940_ (.RESET_B(net277),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0166_),
    .Q(\mydesign.pe_inputs[42] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _5941_ (.RESET_B(net275),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net957),
    .Q(\mydesign.pe_inputs[43] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _5942_ (.RESET_B(net273),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0168_),
    .Q(\mydesign.pe_weights[40] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5943_ (.RESET_B(net271),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0169_),
    .Q(\mydesign.pe_weights[41] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _5944_ (.RESET_B(net269),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0170_),
    .Q(\mydesign.pe_weights[42] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5945_ (.RESET_B(net267),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0171_),
    .Q(\mydesign.pe_weights[43] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _5946_ (.RESET_B(net265),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net740),
    .Q(\mydesign.accum[80] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _5947_ (.RESET_B(net263),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net984),
    .Q(\mydesign.accum[81] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5948_ (.RESET_B(net261),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net962),
    .Q(\mydesign.accum[82] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5949_ (.RESET_B(net259),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0175_),
    .Q(\mydesign.accum[83] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5950_ (.RESET_B(net257),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0176_),
    .Q(\mydesign.accum[84] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5951_ (.RESET_B(net255),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0177_),
    .Q(\mydesign.accum[85] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5952_ (.RESET_B(net253),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0178_),
    .Q(\mydesign.accum[86] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5953_ (.RESET_B(net251),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0179_),
    .Q(\mydesign.accum[87] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _5954_ (.RESET_B(net249),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0180_),
    .Q(\mydesign.pe_inputs[36] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _5955_ (.RESET_B(net247),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0181_),
    .Q(\mydesign.pe_inputs[37] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _5956_ (.RESET_B(net245),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net982),
    .Q(\mydesign.pe_inputs[38] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _5957_ (.RESET_B(net243),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net994),
    .Q(\mydesign.pe_inputs[39] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _5958_ (.RESET_B(net241),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0184_),
    .Q(\mydesign.pe_weights[36] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _5959_ (.RESET_B(net239),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0185_),
    .Q(\mydesign.pe_weights[37] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _5960_ (.RESET_B(net237),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0186_),
    .Q(\mydesign.pe_weights[38] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _5961_ (.RESET_B(net235),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0187_),
    .Q(\mydesign.pe_weights[39] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _5962_ (.RESET_B(net233),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net685),
    .Q(\mydesign.accum[72] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _5963_ (.RESET_B(net231),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net876),
    .Q(\mydesign.accum[73] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _5964_ (.RESET_B(net229),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net883),
    .Q(\mydesign.accum[74] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _5965_ (.RESET_B(net227),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0191_),
    .Q(\mydesign.accum[75] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _5966_ (.RESET_B(net225),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0192_),
    .Q(\mydesign.accum[76] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _5967_ (.RESET_B(net223),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0193_),
    .Q(\mydesign.accum[77] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _5968_ (.RESET_B(net221),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0194_),
    .Q(\mydesign.accum[78] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _5969_ (.RESET_B(net219),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0195_),
    .Q(\mydesign.accum[79] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _5970_ (.RESET_B(net217),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0196_),
    .Q(\mydesign.inputs[3][12] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _5971_ (.RESET_B(net215),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0197_),
    .Q(\mydesign.inputs[3][13] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _5972_ (.RESET_B(net213),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0198_),
    .Q(\mydesign.inputs[3][14] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _5973_ (.RESET_B(net211),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0199_),
    .Q(\mydesign.inputs[3][15] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _5974_ (.RESET_B(net209),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1034),
    .Q(\mydesign.pe_weights[32] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _5975_ (.RESET_B(net207),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0201_),
    .Q(\mydesign.pe_weights[33] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _5976_ (.RESET_B(net205),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0202_),
    .Q(\mydesign.pe_weights[34] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _5977_ (.RESET_B(net203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0203_),
    .Q(\mydesign.pe_weights[35] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _5978_ (.RESET_B(net201),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net691),
    .Q(\mydesign.accum[64] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _5979_ (.RESET_B(net199),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net908),
    .Q(\mydesign.accum[65] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _5980_ (.RESET_B(net197),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net874),
    .Q(\mydesign.accum[66] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _5981_ (.RESET_B(net195),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0207_),
    .Q(\mydesign.accum[67] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _5982_ (.RESET_B(net193),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0208_),
    .Q(\mydesign.accum[68] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _5983_ (.RESET_B(net191),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0209_),
    .Q(\mydesign.accum[69] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _5984_ (.RESET_B(net189),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0210_),
    .Q(\mydesign.accum[70] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _5985_ (.RESET_B(net187),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0211_),
    .Q(\mydesign.accum[71] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _5986_ (.RESET_B(net185),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0212_),
    .Q(\mydesign.pe_inputs[28] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5987_ (.RESET_B(net182),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0213_),
    .Q(\mydesign.pe_inputs[29] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _5988_ (.RESET_B(net178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0214_),
    .Q(\mydesign.pe_inputs[30] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _5989_ (.RESET_B(net170),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0215_),
    .Q(\mydesign.pe_inputs[31] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _5990_ (.RESET_B(net166),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0216_),
    .Q(\mydesign.pe_weights[28] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _5991_ (.RESET_B(net146),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net812),
    .Q(\mydesign.pe_weights[29] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _5992_ (.RESET_B(net142),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net953),
    .Q(\mydesign.pe_weights[30] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5993_ (.RESET_B(net138),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0219_),
    .Q(\mydesign.pe_weights[31] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _5994_ (.RESET_B(net134),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net687),
    .Q(\mydesign.accum[56] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5995_ (.RESET_B(net114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net819),
    .Q(\mydesign.accum[57] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _5996_ (.RESET_B(net110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0222_),
    .Q(\mydesign.accum[58] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _5997_ (.RESET_B(net106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0223_),
    .Q(\mydesign.accum[59] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _5998_ (.RESET_B(net102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0224_),
    .Q(\mydesign.accum[60] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5999_ (.RESET_B(net98),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0225_),
    .Q(\mydesign.accum[61] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6000_ (.RESET_B(net94),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0226_),
    .Q(\mydesign.accum[62] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6001_ (.RESET_B(net90),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0227_),
    .Q(\mydesign.accum[63] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6002_ (.RESET_B(net86),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1023),
    .Q(\mydesign.pe_inputs[24] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6003_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0229_),
    .Q(\mydesign.pe_inputs[25] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6004_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1032),
    .Q(\mydesign.pe_inputs[26] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6005_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net888),
    .Q(\mydesign.pe_inputs[27] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6006_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1014),
    .Q(\mydesign.pe_weights[24] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6007_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net857),
    .Q(\mydesign.pe_weights[25] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6008_ (.RESET_B(net58),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net814),
    .Q(\mydesign.pe_weights[26] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6009_ (.RESET_B(net54),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net790),
    .Q(\mydesign.pe_weights[27] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6010_ (.RESET_B(net50),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net746),
    .Q(\mydesign.accum[48] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6011_ (.RESET_B(net46),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net893),
    .Q(\mydesign.accum[49] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6012_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net901),
    .Q(\mydesign.accum[50] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6013_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0239_),
    .Q(\mydesign.accum[51] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6014_ (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0240_),
    .Q(\mydesign.accum[52] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6015_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0241_),
    .Q(\mydesign.accum[53] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6016_ (.RESET_B(net26),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0242_),
    .Q(\mydesign.accum[54] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6017_ (.RESET_B(net398),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0243_),
    .Q(\mydesign.accum[55] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6018_ (.RESET_B(net394),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0244_),
    .Q(\mydesign.inputs[3][4] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6019_ (.RESET_B(net390),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0245_),
    .Q(\mydesign.inputs[3][5] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6020_ (.RESET_B(net386),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0246_),
    .Q(\mydesign.inputs[3][6] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6021_ (.RESET_B(net382),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0247_),
    .Q(\mydesign.inputs[3][7] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6022_ (.RESET_B(net378),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net846),
    .Q(\mydesign.weights[3][8] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6023_ (.RESET_B(net370),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net860),
    .Q(\mydesign.weights[3][9] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6024_ (.RESET_B(net366),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net855),
    .Q(\mydesign.weights[3][10] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6025_ (.RESET_B(net362),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net822),
    .Q(\mydesign.weights[3][11] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6026_ (.RESET_B(net358),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0252_),
    .Q(\mydesign.pe_inputs[20] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6027_ (.RESET_B(net354),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net850),
    .Q(\mydesign.pe_inputs[21] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6028_ (.RESET_B(net350),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0254_),
    .Q(\mydesign.pe_inputs[22] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6029_ (.RESET_B(net346),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net975),
    .Q(\mydesign.pe_inputs[23] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6030_ (.RESET_B(net342),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0256_),
    .Q(\mydesign.pe_weights[20] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6031_ (.RESET_B(net334),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net863),
    .Q(\mydesign.pe_weights[21] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6032_ (.RESET_B(net330),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net831),
    .Q(\mydesign.pe_weights[22] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6033_ (.RESET_B(net326),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1026),
    .Q(\mydesign.pe_weights[23] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6034_ (.RESET_B(net322),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net665),
    .Q(\mydesign.accum[40] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6035_ (.RESET_B(net318),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net950),
    .Q(\mydesign.accum[41] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6036_ (.RESET_B(net314),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net922),
    .Q(\mydesign.accum[42] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6037_ (.RESET_B(net310),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0263_),
    .Q(\mydesign.accum[43] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6038_ (.RESET_B(net306),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0264_),
    .Q(\mydesign.accum[44] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6039_ (.RESET_B(net302),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0265_),
    .Q(\mydesign.accum[45] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6040_ (.RESET_B(net298),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0266_),
    .Q(\mydesign.accum[46] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6041_ (.RESET_B(net294),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0267_),
    .Q(\mydesign.accum[47] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6042_ (.RESET_B(net290),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net904),
    .Q(\mydesign.pe_weights[16] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6043_ (.RESET_B(net286),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net829),
    .Q(\mydesign.pe_weights[17] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6044_ (.RESET_B(net282),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0270_),
    .Q(\mydesign.pe_weights[18] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6045_ (.RESET_B(net278),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net817),
    .Q(\mydesign.pe_weights[19] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6046_ (.RESET_B(net274),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net735),
    .Q(\mydesign.accum[32] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6047_ (.RESET_B(net270),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net920),
    .Q(\mydesign.accum[33] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6048_ (.RESET_B(net266),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net914),
    .Q(\mydesign.accum[34] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6049_ (.RESET_B(net262),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0275_),
    .Q(\mydesign.accum[35] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6050_ (.RESET_B(net258),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0276_),
    .Q(\mydesign.accum[36] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6051_ (.RESET_B(net254),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0277_),
    .Q(\mydesign.accum[37] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6052_ (.RESET_B(net250),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0278_),
    .Q(\mydesign.accum[38] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _6053_ (.RESET_B(net246),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0279_),
    .Q(\mydesign.accum[39] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6054_ (.RESET_B(net242),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0280_),
    .Q(\mydesign.pe_inputs[12] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6055_ (.RESET_B(net238),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0281_),
    .Q(\mydesign.pe_inputs[13] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6056_ (.RESET_B(net234),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0282_),
    .Q(\mydesign.pe_inputs[14] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6057_ (.RESET_B(net230),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0283_),
    .Q(\mydesign.pe_inputs[15] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6058_ (.RESET_B(net226),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0284_),
    .Q(\mydesign.accum[24] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6059_ (.RESET_B(net222),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net955),
    .Q(\mydesign.accum[25] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6060_ (.RESET_B(net218),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net924),
    .Q(\mydesign.accum[26] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6061_ (.RESET_B(net214),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0287_),
    .Q(\mydesign.accum[27] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6062_ (.RESET_B(net210),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0288_),
    .Q(\mydesign.accum[28] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6063_ (.RESET_B(net206),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0289_),
    .Q(\mydesign.accum[29] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6064_ (.RESET_B(net202),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0290_),
    .Q(\mydesign.accum[30] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6065_ (.RESET_B(net198),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0291_),
    .Q(\mydesign.accum[31] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6066_ (.RESET_B(net194),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net696),
    .Q(\mydesign.weights[2][8] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6067_ (.RESET_B(net192),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net661),
    .Q(\mydesign.weights[2][9] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6068_ (.RESET_B(net190),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net641),
    .Q(\mydesign.weights[2][10] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6069_ (.RESET_B(net188),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net657),
    .Q(\mydesign.weights[2][11] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6070_ (.RESET_B(net186),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1099),
    .Q(\mydesign.pe_inputs[8] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6071_ (.RESET_B(net180),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0297_),
    .Q(\mydesign.pe_inputs[9] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6072_ (.RESET_B(net168),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0298_),
    .Q(\mydesign.pe_inputs[10] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6073_ (.RESET_B(net144),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1001),
    .Q(\mydesign.pe_inputs[11] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6074_ (.RESET_B(net136),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net759),
    .Q(\mydesign.accum[16] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6075_ (.RESET_B(net112),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1030),
    .Q(\mydesign.accum[17] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6076_ (.RESET_B(net104),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1021),
    .Q(\mydesign.accum[18] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6077_ (.RESET_B(net96),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0303_),
    .Q(\mydesign.accum[19] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6078_ (.RESET_B(net88),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0304_),
    .Q(\mydesign.accum[20] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6079_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0305_),
    .Q(\mydesign.accum[21] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6080_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0306_),
    .Q(\mydesign.accum[22] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6081_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0307_),
    .Q(\mydesign.accum[23] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6082_ (.RESET_B(net52),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1066),
    .Q(\mydesign.pe_inputs[4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6083_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net935),
    .Q(\mydesign.pe_inputs[5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6084_ (.RESET_B(net36),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net833),
    .Q(\mydesign.pe_inputs[6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6085_ (.RESET_B(net28),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net947),
    .Q(\mydesign.pe_inputs[7] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6086_ (.RESET_B(net396),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net730),
    .Q(\mydesign.accum[8] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6087_ (.RESET_B(net388),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net929),
    .Q(\mydesign.accum[9] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6088_ (.RESET_B(net380),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1039),
    .Q(\mydesign.accum[10] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6089_ (.RESET_B(net368),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0315_),
    .Q(\mydesign.accum[11] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6090_ (.RESET_B(net360),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0316_),
    .Q(\mydesign.accum[12] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6091_ (.RESET_B(net352),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0317_),
    .Q(\mydesign.accum[13] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6092_ (.RESET_B(net344),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0318_),
    .Q(\mydesign.accum[14] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6093_ (.RESET_B(net332),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1056),
    .Q(\mydesign.accum[15] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6094_ (.RESET_B(net324),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net417),
    .Q(\mydesign.inputs[3][8] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6095_ (.RESET_B(net316),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net659),
    .Q(\mydesign.inputs[3][9] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6096_ (.RESET_B(net308),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net651),
    .Q(\mydesign.inputs[3][10] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6097_ (.RESET_B(net300),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net681),
    .Q(\mydesign.inputs[3][11] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _6098_ (.RESET_B(net292),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net750),
    .Q(\mydesign.accum[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6099_ (.RESET_B(net284),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1058),
    .Q(\mydesign.accum[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6100_ (.RESET_B(net276),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1041),
    .Q(\mydesign.accum[2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6101_ (.RESET_B(net268),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0327_),
    .Q(\mydesign.accum[3] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6102_ (.RESET_B(net260),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0328_),
    .Q(\mydesign.accum[4] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6103_ (.RESET_B(net252),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0329_),
    .Q(\mydesign.accum[5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6104_ (.RESET_B(net244),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0330_),
    .Q(\mydesign.accum[6] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6105_ (.RESET_B(net236),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net410),
    .Q(\mydesign.accum[7] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6106_ (.RESET_B(net228),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0332_),
    .Q(\mydesign.weights[1][16] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6107_ (.RESET_B(net224),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0333_),
    .Q(\mydesign.weights[1][17] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6108_ (.RESET_B(net220),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0334_),
    .Q(\mydesign.weights[1][18] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6109_ (.RESET_B(net216),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0335_),
    .Q(\mydesign.weights[1][19] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6110_ (.RESET_B(net212),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0336_),
    .Q(\mydesign.out[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _6111_ (.RESET_B(net204),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0337_),
    .Q(\mydesign.out[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6112_ (.RESET_B(net196),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0338_),
    .Q(\mydesign.out[2] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6113_ (.RESET_B(net176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1104),
    .Q(\mydesign.out[3] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6114_ (.RESET_B(net140),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net726),
    .Q(\mydesign.weights[3][0] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6115_ (.RESET_B(net132),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net718),
    .Q(\mydesign.weights[3][1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6116_ (.RESET_B(net108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net706),
    .Q(\mydesign.weights[3][2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6117_ (.RESET_B(net100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net732),
    .Q(\mydesign.weights[3][3] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6118_ (.RESET_B(net92),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0344_),
    .Q(\mydesign.weights[1][8] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6119_ (.RESET_B(net84),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0345_),
    .Q(\mydesign.weights[1][9] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6120_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0346_),
    .Q(\mydesign.weights[1][10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6121_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0347_),
    .Q(\mydesign.weights[1][11] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6122_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0348_),
    .Q(\mydesign.weights[1][12] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6123_ (.RESET_B(net48),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0349_),
    .Q(\mydesign.weights[1][13] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6124_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0350_),
    .Q(\mydesign.weights[1][14] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6125_ (.RESET_B(net32),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0351_),
    .Q(\mydesign.weights[1][15] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6126_ (.RESET_B(net24),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net724),
    .Q(\mydesign.weights[0][24] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6127_ (.RESET_B(net392),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0353_),
    .Q(\mydesign.weights[0][25] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6128_ (.RESET_B(net384),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0354_),
    .Q(\mydesign.weights[0][26] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6129_ (.RESET_B(net372),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net715),
    .Q(\mydesign.weights[0][27] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6130_ (.RESET_B(net364),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0356_),
    .Q(\mydesign.weights[0][20] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6131_ (.RESET_B(net356),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0357_),
    .Q(\mydesign.weights[0][21] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6132_ (.RESET_B(net348),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0358_),
    .Q(\mydesign.weights[0][22] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6133_ (.RESET_B(net336),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0359_),
    .Q(\mydesign.weights[0][23] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6134_ (.RESET_B(net328),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0360_),
    .Q(\mydesign.weights[0][16] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6135_ (.RESET_B(net320),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0361_),
    .Q(\mydesign.weights[0][17] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6136_ (.RESET_B(net312),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0362_),
    .Q(\mydesign.weights[0][18] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6137_ (.RESET_B(net304),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0363_),
    .Q(\mydesign.weights[0][19] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6138_ (.RESET_B(net296),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net987),
    .Q(\mydesign.weights[3][12] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6139_ (.RESET_B(net280),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net825),
    .Q(\mydesign.weights[3][13] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6140_ (.RESET_B(net264),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net932),
    .Q(\mydesign.weights[3][14] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6141_ (.RESET_B(net248),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net871),
    .Q(\mydesign.weights[3][15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6142_ (.RESET_B(net232),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0368_),
    .Q(\mydesign.weights[0][12] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6143_ (.RESET_B(net208),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0369_),
    .Q(\mydesign.weights[0][13] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6144_ (.RESET_B(net200),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0370_),
    .Q(\mydesign.weights[0][14] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6145_ (.RESET_B(net184),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0371_),
    .Q(\mydesign.weights[0][15] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6146_ (.RESET_B(net164),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0372_),
    .Q(\mydesign.weights[1][20] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6147_ (.RESET_B(net288),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0373_),
    .Q(\mydesign.weights[1][21] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6148_ (.RESET_B(net272),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0374_),
    .Q(\mydesign.weights[1][22] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6149_ (.RESET_B(net256),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0375_),
    .Q(\mydesign.weights[1][23] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_tiehi _6126__24 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net24));
 sg13g2_tiehi _5874__25 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net25));
 sg13g2_tiehi _6016__26 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net26));
 sg13g2_tiehi _5873__27 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net27));
 sg13g2_tiehi _6085__28 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net28));
 sg13g2_tiehi _5872__29 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net29));
 sg13g2_tiehi _6015__30 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net30));
 sg13g2_tiehi _5871__31 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net31));
 sg13g2_tiehi _6125__32 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net32));
 sg13g2_tiehi _5870__33 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net33));
 sg13g2_tiehi _6014__34 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net34));
 sg13g2_tiehi _5869__35 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net35));
 sg13g2_tiehi _6084__36 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net36));
 sg13g2_tiehi _5868__37 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net37));
 sg13g2_tiehi _6013__38 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net38));
 sg13g2_tiehi _5867__39 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_tiehi _6124__40 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_tiehi _5866__41 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net41));
 sg13g2_tiehi _6012__42 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net42));
 sg13g2_tiehi _5865__43 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net43));
 sg13g2_tiehi _6083__44 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net44));
 sg13g2_tiehi _5864__45 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net45));
 sg13g2_tiehi _6011__46 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net46));
 sg13g2_tiehi _5863__47 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net47));
 sg13g2_tiehi _6123__48 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net48));
 sg13g2_tiehi _5862__49 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net49));
 sg13g2_tiehi _6010__50 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net50));
 sg13g2_tiehi _5861__51 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net51));
 sg13g2_tiehi _6082__52 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net52));
 sg13g2_tiehi _5860__53 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net53));
 sg13g2_tiehi _6009__54 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net54));
 sg13g2_tiehi _5859__55 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net55));
 sg13g2_tiehi _6122__56 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net56));
 sg13g2_tiehi _5858__57 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net57));
 sg13g2_tiehi _6008__58 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net58));
 sg13g2_tiehi _5857__59 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net59));
 sg13g2_tiehi _6081__60 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net60));
 sg13g2_tiehi _5856__61 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net61));
 sg13g2_tiehi _6007__62 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net62));
 sg13g2_tiehi _5855__63 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net63));
 sg13g2_tiehi _6121__64 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net64));
 sg13g2_tiehi _5854__65 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net65));
 sg13g2_tiehi _5853__66 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net66));
 sg13g2_tiehi _5852__67 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net67));
 sg13g2_tiehi _5851__68 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net68));
 sg13g2_tiehi _5850__69 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net69));
 sg13g2_tiehi _6006__70 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net70));
 sg13g2_tiehi _5849__71 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net71));
 sg13g2_tiehi _6080__72 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net72));
 sg13g2_tiehi _5848__73 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net73));
 sg13g2_tiehi _6005__74 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net74));
 sg13g2_tiehi _5847__75 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net75));
 sg13g2_tiehi _6120__76 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net76));
 sg13g2_tiehi _5846__77 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net77));
 sg13g2_tiehi _6004__78 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net78));
 sg13g2_tiehi _5845__79 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net79));
 sg13g2_tiehi _6079__80 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net80));
 sg13g2_tiehi _5844__81 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net81));
 sg13g2_tiehi _6003__82 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net82));
 sg13g2_tiehi _5843__83 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net83));
 sg13g2_tiehi _6119__84 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net84));
 sg13g2_tiehi _5842__85 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net85));
 sg13g2_tiehi _6002__86 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net86));
 sg13g2_tiehi _5841__87 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net87));
 sg13g2_tiehi _6078__88 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net88));
 sg13g2_tiehi _5840__89 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net89));
 sg13g2_tiehi _6001__90 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net90));
 sg13g2_tiehi _5839__91 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net91));
 sg13g2_tiehi _6118__92 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net92));
 sg13g2_tiehi _5838__93 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net93));
 sg13g2_tiehi _6000__94 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net94));
 sg13g2_tiehi _5837__95 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net95));
 sg13g2_tiehi _6077__96 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net96));
 sg13g2_tiehi _5836__97 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net97));
 sg13g2_tiehi _5999__98 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net98));
 sg13g2_tiehi _5835__99 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net99));
 sg13g2_tiehi _6117__100 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net100));
 sg13g2_tiehi _5834__101 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net101));
 sg13g2_tiehi _5998__102 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net102));
 sg13g2_tiehi _5833__103 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net103));
 sg13g2_tiehi _6076__104 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net104));
 sg13g2_tiehi _5832__105 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net105));
 sg13g2_tiehi _5997__106 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net106));
 sg13g2_tiehi _5831__107 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net107));
 sg13g2_tiehi _6116__108 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net108));
 sg13g2_tiehi _5830__109 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net109));
 sg13g2_tiehi _5996__110 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net110));
 sg13g2_tiehi _5829__111 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net111));
 sg13g2_tiehi _6075__112 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net112));
 sg13g2_tiehi _5828__113 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net113));
 sg13g2_tiehi _5995__114 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net114));
 sg13g2_tiehi _5827__115 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net115));
 sg13g2_tiehi _5826__116 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net116));
 sg13g2_tiehi _5825__117 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net117));
 sg13g2_tiehi _5824__118 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net118));
 sg13g2_tiehi _5823__119 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net119));
 sg13g2_tiehi _5822__120 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net120));
 sg13g2_tiehi _5821__121 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net121));
 sg13g2_tiehi _5820__122 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net122));
 sg13g2_tiehi _5819__123 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net123));
 sg13g2_tiehi _5818__124 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net124));
 sg13g2_tiehi _5817__125 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net125));
 sg13g2_tiehi _5816__126 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net126));
 sg13g2_tiehi _5815__127 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net127));
 sg13g2_tiehi _5814__128 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net128));
 sg13g2_tiehi _5813__129 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net129));
 sg13g2_tiehi _5812__130 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net130));
 sg13g2_tiehi _5811__131 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net131));
 sg13g2_tiehi _6115__132 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net132));
 sg13g2_tiehi _5810__133 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net133));
 sg13g2_tiehi _5994__134 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net134));
 sg13g2_tiehi _5809__135 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net135));
 sg13g2_tiehi _6074__136 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net136));
 sg13g2_tiehi _5808__137 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net137));
 sg13g2_tiehi _5993__138 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net138));
 sg13g2_tiehi _5807__139 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net139));
 sg13g2_tiehi _6114__140 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net140));
 sg13g2_tiehi _5806__141 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net141));
 sg13g2_tiehi _5992__142 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net142));
 sg13g2_tiehi _5805__143 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net143));
 sg13g2_tiehi _6073__144 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net144));
 sg13g2_tiehi _5804__145 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net145));
 sg13g2_tiehi _5991__146 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net146));
 sg13g2_tiehi _5803__147 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net147));
 sg13g2_tiehi _5802__148 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net148));
 sg13g2_tiehi _5801__149 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net149));
 sg13g2_tiehi _5800__150 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net150));
 sg13g2_tiehi _5799__151 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net151));
 sg13g2_tiehi _5798__152 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net152));
 sg13g2_tiehi _5797__153 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net153));
 sg13g2_tiehi _5796__154 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net154));
 sg13g2_tiehi _5795__155 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net155));
 sg13g2_tiehi _5794__156 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net156));
 sg13g2_tiehi _5793__157 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net157));
 sg13g2_tiehi _5792__158 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net158));
 sg13g2_tiehi _5791__159 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net159));
 sg13g2_tiehi _5790__160 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net160));
 sg13g2_tiehi _5789__161 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net161));
 sg13g2_tiehi _5788__162 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net162));
 sg13g2_tiehi _5787__163 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net163));
 sg13g2_tiehi _6146__164 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net164));
 sg13g2_tiehi _5786__165 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net165));
 sg13g2_tiehi _5990__166 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net166));
 sg13g2_tiehi _5785__167 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net167));
 sg13g2_tiehi _6072__168 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net168));
 sg13g2_tiehi _5784__169 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net169));
 sg13g2_tiehi _5989__170 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net170));
 sg13g2_tiehi _5783__171 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net171));
 sg13g2_tiehi _5782__172 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net172));
 sg13g2_tiehi _5781__173 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net173));
 sg13g2_tiehi _5780__174 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net174));
 sg13g2_tiehi _5779__175 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net175));
 sg13g2_tiehi _6113__176 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net176));
 sg13g2_tiehi _5778__177 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net177));
 sg13g2_tiehi _5988__178 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net178));
 sg13g2_tiehi _5777__179 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net179));
 sg13g2_tiehi _6071__180 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net180));
 sg13g2_tiehi _5776__181 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net181));
 sg13g2_tiehi _5987__182 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net182));
 sg13g2_tiehi _5775__183 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net183));
 sg13g2_tiehi _6145__184 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net184));
 sg13g2_tiehi _5986__185 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net185));
 sg13g2_tiehi _6070__186 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net186));
 sg13g2_tiehi _5985__187 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net187));
 sg13g2_tiehi _6069__188 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net188));
 sg13g2_tiehi _5984__189 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net189));
 sg13g2_tiehi _6068__190 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net190));
 sg13g2_tiehi _5983__191 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net191));
 sg13g2_tiehi _6067__192 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net192));
 sg13g2_tiehi _5982__193 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net193));
 sg13g2_tiehi _6066__194 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net194));
 sg13g2_tiehi _5981__195 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net195));
 sg13g2_tiehi _6112__196 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net196));
 sg13g2_tiehi _5980__197 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net197));
 sg13g2_tiehi _6065__198 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net198));
 sg13g2_tiehi _5979__199 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net199));
 sg13g2_tiehi _6144__200 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net200));
 sg13g2_tiehi _5978__201 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net201));
 sg13g2_tiehi _6064__202 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net202));
 sg13g2_tiehi _5977__203 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net203));
 sg13g2_tiehi _6111__204 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net204));
 sg13g2_tiehi _5976__205 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net205));
 sg13g2_tiehi _6063__206 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net206));
 sg13g2_tiehi _5975__207 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net207));
 sg13g2_tiehi _6143__208 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net208));
 sg13g2_tiehi _5974__209 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net209));
 sg13g2_tiehi _6062__210 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net210));
 sg13g2_tiehi _5973__211 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net211));
 sg13g2_tiehi _6110__212 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net212));
 sg13g2_tiehi _5972__213 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net213));
 sg13g2_tiehi _6061__214 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net214));
 sg13g2_tiehi _5971__215 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net215));
 sg13g2_tiehi _6109__216 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net216));
 sg13g2_tiehi _5970__217 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net217));
 sg13g2_tiehi _6060__218 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net218));
 sg13g2_tiehi _5969__219 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net219));
 sg13g2_tiehi _6108__220 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net220));
 sg13g2_tiehi _5968__221 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net221));
 sg13g2_tiehi _6059__222 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net222));
 sg13g2_tiehi _5967__223 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net223));
 sg13g2_tiehi _6107__224 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net224));
 sg13g2_tiehi _5966__225 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net225));
 sg13g2_tiehi _6058__226 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net226));
 sg13g2_tiehi _5965__227 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net227));
 sg13g2_tiehi _6106__228 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net228));
 sg13g2_tiehi _5964__229 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net229));
 sg13g2_tiehi _6057__230 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net230));
 sg13g2_tiehi _5963__231 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net231));
 sg13g2_tiehi _6142__232 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net232));
 sg13g2_tiehi _5962__233 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net233));
 sg13g2_tiehi _6056__234 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net234));
 sg13g2_tiehi _5961__235 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net235));
 sg13g2_tiehi _6105__236 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net236));
 sg13g2_tiehi _5960__237 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net237));
 sg13g2_tiehi _6055__238 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net238));
 sg13g2_tiehi _5959__239 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net239));
 sg13g2_tiehi _5774__240 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net240));
 sg13g2_tiehi _5958__241 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net241));
 sg13g2_tiehi _6054__242 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net242));
 sg13g2_tiehi _5957__243 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net243));
 sg13g2_tiehi _6104__244 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net244));
 sg13g2_tiehi _5956__245 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net245));
 sg13g2_tiehi _6053__246 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net246));
 sg13g2_tiehi _5955__247 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net247));
 sg13g2_tiehi _6141__248 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net248));
 sg13g2_tiehi _5954__249 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net249));
 sg13g2_tiehi _6052__250 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net250));
 sg13g2_tiehi _5953__251 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net251));
 sg13g2_tiehi _6103__252 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net252));
 sg13g2_tiehi _5952__253 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net253));
 sg13g2_tiehi _6051__254 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net254));
 sg13g2_tiehi _5951__255 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net255));
 sg13g2_tiehi _6149__256 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net256));
 sg13g2_tiehi _5950__257 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net257));
 sg13g2_tiehi _6050__258 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net258));
 sg13g2_tiehi _5949__259 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net259));
 sg13g2_tiehi _6102__260 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net260));
 sg13g2_tiehi _5948__261 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net261));
 sg13g2_tiehi _6049__262 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net262));
 sg13g2_tiehi _5947__263 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net263));
 sg13g2_tiehi _6140__264 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net264));
 sg13g2_tiehi _5946__265 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net265));
 sg13g2_tiehi _6048__266 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net266));
 sg13g2_tiehi _5945__267 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net267));
 sg13g2_tiehi _6101__268 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net268));
 sg13g2_tiehi _5944__269 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net269));
 sg13g2_tiehi _6047__270 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net270));
 sg13g2_tiehi _5943__271 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net271));
 sg13g2_tiehi _6148__272 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net272));
 sg13g2_tiehi _5942__273 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net273));
 sg13g2_tiehi _6046__274 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net274));
 sg13g2_tiehi _5941__275 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net275));
 sg13g2_tiehi _6100__276 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net276));
 sg13g2_tiehi _5940__277 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net277));
 sg13g2_tiehi _6045__278 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net278));
 sg13g2_tiehi _5939__279 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net279));
 sg13g2_tiehi _6139__280 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net280));
 sg13g2_tiehi _5938__281 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net281));
 sg13g2_tiehi _6044__282 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net282));
 sg13g2_tiehi _5937__283 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net283));
 sg13g2_tiehi _6099__284 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net284));
 sg13g2_tiehi _5936__285 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net285));
 sg13g2_tiehi _6043__286 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net286));
 sg13g2_tiehi _5935__287 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net287));
 sg13g2_tiehi _6147__288 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net288));
 sg13g2_tiehi _5934__289 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net289));
 sg13g2_tiehi _6042__290 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net290));
 sg13g2_tiehi _5933__291 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net291));
 sg13g2_tiehi _6098__292 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net292));
 sg13g2_tiehi _5932__293 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net293));
 sg13g2_tiehi _6041__294 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net294));
 sg13g2_tiehi _5931__295 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net295));
 sg13g2_tiehi _6138__296 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net296));
 sg13g2_tiehi _5930__297 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net297));
 sg13g2_tiehi _6040__298 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net298));
 sg13g2_tiehi _5929__299 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net299));
 sg13g2_tiehi _6097__300 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net300));
 sg13g2_tiehi _5928__301 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net301));
 sg13g2_tiehi _6039__302 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net302));
 sg13g2_tiehi _5927__303 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net303));
 sg13g2_tiehi _6137__304 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net304));
 sg13g2_tiehi _5926__305 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net305));
 sg13g2_tiehi _6038__306 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net306));
 sg13g2_tiehi _5925__307 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net307));
 sg13g2_tiehi _6096__308 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net308));
 sg13g2_tiehi _5924__309 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net309));
 sg13g2_tiehi _6037__310 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net310));
 sg13g2_tiehi _5923__311 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net311));
 sg13g2_tiehi _6136__312 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net312));
 sg13g2_tiehi _5922__313 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net313));
 sg13g2_tiehi _6036__314 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net314));
 sg13g2_tiehi _5921__315 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net315));
 sg13g2_tiehi _6095__316 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net316));
 sg13g2_tiehi _5920__317 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net317));
 sg13g2_tiehi _6035__318 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net318));
 sg13g2_tiehi _5919__319 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net319));
 sg13g2_tiehi _6135__320 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net320));
 sg13g2_tiehi _5918__321 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net321));
 sg13g2_tiehi _6034__322 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net322));
 sg13g2_tiehi _5917__323 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net323));
 sg13g2_tiehi _6094__324 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net324));
 sg13g2_tiehi _5916__325 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net325));
 sg13g2_tiehi _6033__326 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net326));
 sg13g2_tiehi _5915__327 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net327));
 sg13g2_tiehi _6134__328 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net328));
 sg13g2_tiehi _5914__329 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net329));
 sg13g2_tiehi _6032__330 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net330));
 sg13g2_tiehi _5913__331 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net331));
 sg13g2_tiehi _6093__332 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net332));
 sg13g2_tiehi _5912__333 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net333));
 sg13g2_tiehi _6031__334 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net334));
 sg13g2_tiehi _5911__335 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net335));
 sg13g2_tiehi _6133__336 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net336));
 sg13g2_tiehi _5910__337 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net337));
 sg13g2_tiehi _5909__338 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net338));
 sg13g2_tiehi _5908__339 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net339));
 sg13g2_tiehi _5907__340 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net340));
 sg13g2_tiehi _5906__341 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net341));
 sg13g2_tiehi _6030__342 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net342));
 sg13g2_tiehi _5905__343 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net343));
 sg13g2_tiehi _6092__344 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net344));
 sg13g2_tiehi _5904__345 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net345));
 sg13g2_tiehi _6029__346 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net346));
 sg13g2_tiehi _5903__347 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net347));
 sg13g2_tiehi _6132__348 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net348));
 sg13g2_tiehi _5902__349 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net349));
 sg13g2_tiehi _6028__350 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net350));
 sg13g2_tiehi _5901__351 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net351));
 sg13g2_tiehi _6091__352 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net352));
 sg13g2_tiehi _5900__353 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net353));
 sg13g2_tiehi _6027__354 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net354));
 sg13g2_tiehi _5899__355 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net355));
 sg13g2_tiehi _6131__356 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net356));
 sg13g2_tiehi _5898__357 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net357));
 sg13g2_tiehi _6026__358 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net358));
 sg13g2_tiehi _5897__359 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net359));
 sg13g2_tiehi _6090__360 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net360));
 sg13g2_tiehi _5896__361 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net361));
 sg13g2_tiehi _6025__362 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net362));
 sg13g2_tiehi _5895__363 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net363));
 sg13g2_tiehi _6130__364 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net364));
 sg13g2_tiehi _5894__365 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net365));
 sg13g2_tiehi _6024__366 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net366));
 sg13g2_tiehi _5893__367 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net367));
 sg13g2_tiehi _6089__368 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net368));
 sg13g2_tiehi _5892__369 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net369));
 sg13g2_tiehi _6023__370 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net370));
 sg13g2_tiehi _5891__371 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net371));
 sg13g2_tiehi _6129__372 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net372));
 sg13g2_tiehi _5890__373 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net373));
 sg13g2_tiehi _5889__374 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net374));
 sg13g2_tiehi _5888__375 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net375));
 sg13g2_tiehi _5887__376 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net376));
 sg13g2_tiehi _5886__377 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net377));
 sg13g2_tiehi _6022__378 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net378));
 sg13g2_tiehi _5885__379 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net379));
 sg13g2_tiehi _6088__380 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net380));
 sg13g2_tiehi _5884__381 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net381));
 sg13g2_tiehi _6021__382 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net382));
 sg13g2_tiehi _5883__383 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net383));
 sg13g2_tiehi _6128__384 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net384));
 sg13g2_tiehi _5882__385 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net385));
 sg13g2_tiehi _6020__386 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net386));
 sg13g2_tiehi _5881__387 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net387));
 sg13g2_tiehi _6087__388 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net388));
 sg13g2_tiehi _5880__389 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net389));
 sg13g2_tiehi _6019__390 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net390));
 sg13g2_tiehi _5879__391 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net391));
 sg13g2_tiehi _6127__392 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net392));
 sg13g2_tiehi _5878__393 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net393));
 sg13g2_tiehi _6018__394 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net394));
 sg13g2_tiehi _5877__395 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net395));
 sg13g2_tiehi _6086__396 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net396));
 sg13g2_tiehi _5876__397 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net397));
 sg13g2_tiehi _6017__398 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net398));
 sg13g2_tiehi heichips25_systolicArrayTop_399 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net399));
 sg13g2_tiehi heichips25_systolicArrayTop_400 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net400));
 sg13g2_tiehi heichips25_systolicArrayTop_401 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net401));
 sg13g2_tiehi heichips25_systolicArrayTop_402 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net402));
 sg13g2_tiehi heichips25_systolicArrayTop_403 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net403));
 sg13g2_tiehi heichips25_systolicArrayTop_404 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net404));
 sg13g2_tiehi heichips25_systolicArrayTop_405 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net405));
 sg13g2_tiehi heichips25_systolicArrayTop_406 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net406));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_systolicArrayTop_17 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net17));
 sg13g2_tielo heichips25_systolicArrayTop_18 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net18));
 sg13g2_tielo heichips25_systolicArrayTop_19 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net19));
 sg13g2_tielo heichips25_systolicArrayTop_20 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net20));
 sg13g2_tielo heichips25_systolicArrayTop_21 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net21));
 sg13g2_tielo heichips25_systolicArrayTop_22 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net22));
 sg13g2_tiehi _5875__23 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net23));
 sg13g2_buf_1 _6541_ (.A(\mydesign.valid_out ),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout428 (.A(_0933_),
    .X(net428),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout429 (.A(_2692_),
    .X(net429),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout430 (.A(net431),
    .X(net430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout431 (.A(_2697_),
    .X(net431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout432 (.A(_2608_),
    .X(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout433 (.A(net435),
    .X(net433),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout434 (.A(net435),
    .X(net434),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout435 (.A(net439),
    .X(net435),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout436 (.A(net437),
    .X(net436),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout437 (.A(net438),
    .X(net437),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout438 (.A(net439),
    .X(net438),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout439 (.A(net453),
    .X(net439),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout440 (.A(net441),
    .X(net440),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout441 (.A(net453),
    .X(net441),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout442 (.A(net446),
    .X(net442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout443 (.A(net446),
    .X(net443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout444 (.A(net445),
    .X(net444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout445 (.A(net446),
    .X(net445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout446 (.A(net453),
    .X(net446),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout447 (.A(net452),
    .X(net447),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout448 (.A(net452),
    .X(net448),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout449 (.A(net450),
    .X(net449),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout450 (.A(net451),
    .X(net450),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout451 (.A(net452),
    .X(net451),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout452 (.A(net453),
    .X(net452),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout453 (.A(_2601_),
    .X(net453),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout454 (.A(_2596_),
    .X(net454),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout455 (.A(_0498_),
    .X(net455),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout456 (.A(_0407_),
    .X(net456),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout457 (.A(net458),
    .X(net457),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout458 (.A(_0403_),
    .X(net458),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout459 (.A(_0396_),
    .X(net459),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout460 (.A(_0396_),
    .X(net460),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout461 (.A(_0390_),
    .X(net461),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout462 (.A(_2661_),
    .X(net462),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout463 (.A(_2661_),
    .X(net463),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout464 (.A(net466),
    .X(net464),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout465 (.A(net466),
    .X(net465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout466 (.A(net483),
    .X(net466),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout467 (.A(net469),
    .X(net467),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout468 (.A(net469),
    .X(net468),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout469 (.A(net483),
    .X(net469),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout470 (.A(net472),
    .X(net470),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout471 (.A(net472),
    .X(net471),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout472 (.A(net483),
    .X(net472),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout473 (.A(net474),
    .X(net473),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout474 (.A(net478),
    .X(net474),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout475 (.A(net477),
    .X(net475),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout476 (.A(net477),
    .X(net476),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout477 (.A(net478),
    .X(net477),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout478 (.A(net483),
    .X(net478),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout479 (.A(net480),
    .X(net479),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout480 (.A(net482),
    .X(net480),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout481 (.A(net482),
    .X(net481),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout482 (.A(net483),
    .X(net482),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout483 (.A(_2660_),
    .X(net483),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout484 (.A(net485),
    .X(net484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout485 (.A(_2602_),
    .X(net485),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout486 (.A(net490),
    .X(net486),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout487 (.A(net490),
    .X(net487),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout488 (.A(net490),
    .X(net488),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout489 (.A(net490),
    .X(net489),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout490 (.A(_2602_),
    .X(net490),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout491 (.A(net494),
    .X(net491),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout492 (.A(net494),
    .X(net492),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout493 (.A(net494),
    .X(net493),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout494 (.A(_2602_),
    .X(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout495 (.A(net496),
    .X(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout496 (.A(_2595_),
    .X(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout497 (.A(_2587_),
    .X(net497),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout498 (.A(_2587_),
    .X(net498),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout499 (.A(_2516_),
    .X(net499),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout500 (.A(_2516_),
    .X(net500),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout501 (.A(net503),
    .X(net501),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout502 (.A(net503),
    .X(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout503 (.A(_2516_),
    .X(net503),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout504 (.A(net510),
    .X(net504),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout505 (.A(net510),
    .X(net505),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout506 (.A(net507),
    .X(net506),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout507 (.A(net510),
    .X(net507),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout508 (.A(net509),
    .X(net508),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout509 (.A(net510),
    .X(net509),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout510 (.A(net1103),
    .X(net510),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout511 (.A(net518),
    .X(net511),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout512 (.A(net518),
    .X(net512),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout513 (.A(net514),
    .X(net513),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout514 (.A(net517),
    .X(net514),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout515 (.A(net516),
    .X(net515),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout516 (.A(net517),
    .X(net516),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout517 (.A(net518),
    .X(net517),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout518 (.A(net1105),
    .X(net518),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout519 (.A(\mydesign.pe_inputs[7] ),
    .X(net519),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout520 (.A(\mydesign.pe_inputs[11] ),
    .X(net520),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout521 (.A(\mydesign.pe_inputs[8] ),
    .X(net521),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout522 (.A(net1098),
    .X(net522),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout523 (.A(net524),
    .X(net523),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout524 (.A(net903),
    .X(net524),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout525 (.A(\mydesign.pe_weights[22] ),
    .X(net525),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout526 (.A(net1097),
    .X(net526),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout527 (.A(\mydesign.pe_weights[27] ),
    .X(net527),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout528 (.A(net1022),
    .X(net528),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout529 (.A(net1094),
    .X(net529),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout530 (.A(net938),
    .X(net530),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout531 (.A(net1101),
    .X(net531),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout532 (.A(net1095),
    .X(net532),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout533 (.A(net789),
    .X(net533),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout534 (.A(net1050),
    .X(net534),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout535 (.A(net927),
    .X(net535),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout536 (.A(net1100),
    .X(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout537 (.A(net1067),
    .X(net537),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout538 (.A(net1092),
    .X(net538),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout539 (.A(net1096),
    .X(net539),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout540 (.A(net1102),
    .X(net540),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout541 (.A(net543),
    .X(net541),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout542 (.A(net543),
    .X(net542),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout543 (.A(net1083),
    .X(net543),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout544 (.A(net545),
    .X(net544),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout545 (.A(net546),
    .X(net545),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout546 (.A(net1088),
    .X(net546),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout547 (.A(net548),
    .X(net547),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout548 (.A(net553),
    .X(net548),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout549 (.A(net552),
    .X(net549),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout550 (.A(net552),
    .X(net550),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout551 (.A(net552),
    .X(net551),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout552 (.A(net553),
    .X(net552),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout553 (.A(\mydesign.cp[0] ),
    .X(net553),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout554 (.A(net556),
    .X(net554),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout555 (.A(net556),
    .X(net555),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout556 (.A(net557),
    .X(net556),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout557 (.A(\mydesign.cp[0] ),
    .X(net557),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout558 (.A(net562),
    .X(net558),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout559 (.A(net562),
    .X(net559),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout560 (.A(net562),
    .X(net560),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout561 (.A(net562),
    .X(net561),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout562 (.A(net595),
    .X(net562),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout563 (.A(net595),
    .X(net563),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout564 (.A(net565),
    .X(net564),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout565 (.A(net566),
    .X(net565),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout566 (.A(net571),
    .X(net566),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout567 (.A(net569),
    .X(net567),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout568 (.A(net569),
    .X(net568),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout569 (.A(net571),
    .X(net569),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout570 (.A(net571),
    .X(net570),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout571 (.A(net595),
    .X(net571),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout572 (.A(net573),
    .X(net572),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout573 (.A(net576),
    .X(net573),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout574 (.A(net576),
    .X(net574),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout575 (.A(net576),
    .X(net575),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout576 (.A(net594),
    .X(net576),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout577 (.A(net578),
    .X(net577),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout578 (.A(net581),
    .X(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout579 (.A(net580),
    .X(net579),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout581 (.A(net594),
    .X(net581),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout582 (.A(net583),
    .X(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout583 (.A(net594),
    .X(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout584 (.A(net585),
    .X(net584),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout585 (.A(net589),
    .X(net585),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout586 (.A(net587),
    .X(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout587 (.A(net588),
    .X(net587),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout588 (.A(net589),
    .X(net588),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout589 (.A(net594),
    .X(net589),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout590 (.A(net591),
    .X(net590),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout591 (.A(net593),
    .X(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout592 (.A(net593),
    .X(net592),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout593 (.A(net594),
    .X(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout594 (.A(net595),
    .X(net594),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout595 (.A(net867),
    .X(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout596 (.A(net1093),
    .X(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout597 (.A(_2631_),
    .X(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout598 (.A(_2631_),
    .X(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout599 (.A(_2629_),
    .X(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout600 (.A(_2629_),
    .X(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout601 (.A(_2627_),
    .X(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout602 (.A(_2627_),
    .X(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout603 (.A(_2625_),
    .X(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout604 (.A(_2625_),
    .X(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout605 (.A(_2617_),
    .X(net605),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout606 (.A(_2617_),
    .X(net606),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout607 (.A(net608),
    .X(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout608 (.A(net609),
    .X(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout609 (.A(_2590_),
    .X(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout610 (.A(net611),
    .X(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout611 (.A(ui_in[4]),
    .X(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout612 (.A(net613),
    .X(net612),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout613 (.A(net619),
    .X(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout614 (.A(net615),
    .X(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout615 (.A(net619),
    .X(net615),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout616 (.A(net617),
    .X(net616),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout617 (.A(net619),
    .X(net617),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout618 (.A(net619),
    .X(net618),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout619 (.A(net640),
    .X(net619),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout620 (.A(net621),
    .X(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout621 (.A(net640),
    .X(net621),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout622 (.A(net623),
    .X(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout623 (.A(net627),
    .X(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout624 (.A(net627),
    .X(net624),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout625 (.A(net626),
    .X(net625),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout626 (.A(net627),
    .X(net626),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout627 (.A(net640),
    .X(net627),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout628 (.A(net632),
    .X(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout629 (.A(net632),
    .X(net629),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout630 (.A(net632),
    .X(net630),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout631 (.A(net632),
    .X(net631),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout632 (.A(net639),
    .X(net632),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout633 (.A(net636),
    .X(net633),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout634 (.A(net636),
    .X(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout635 (.A(net636),
    .X(net635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout636 (.A(net639),
    .X(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout637 (.A(net639),
    .X(net637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout638 (.A(net639),
    .X(net638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout639 (.A(net640),
    .X(net639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout640 (.A(rst_n),
    .X(net640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input5 (.A(ui_in[5]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input6 (.A(ui_in[6]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_systolicArrayTop_16 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net16));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_14_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_30_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_39_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_40_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_41_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_42_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_43_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_44_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_45_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_46_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_47_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_48_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_49_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload0 (.A(clknet_3_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload1 (.A(clknet_3_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload2 (.A(clknet_3_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload3 (.A(clknet_3_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload4 (.A(clknet_3_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload5 (.A(clknet_3_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_49_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload10 (.A(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload11 (.VDD(VPWR),
    .A(clknet_leaf_39_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload12 (.VDD(VPWR),
    .A(clknet_leaf_41_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload14 (.VDD(VPWR),
    .A(clknet_leaf_34_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload15 (.VDD(VPWR),
    .A(clknet_leaf_37_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload17 (.A(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload18 (.VDD(VPWR),
    .A(clknet_leaf_33_clk),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mydesign.cp2[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0067_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mydesign.accum[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0331_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mydesign.weights[3][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0112_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mydesign.inputs[2][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mydesign.inputs[2][12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0076_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mydesign.inputs[3][8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0320_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mydesign.inputs[2][14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0078_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mydesign.inputs[2][9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0014_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mydesign.inputs[3][14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mydesign.inputs[2][8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0013_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold19 (.A(\mydesign.inputs[2][13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0077_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mydesign.weights[2][10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0294_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mydesign.inputs[2][11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0016_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold25 (.A(\mydesign.inputs[3][13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mydesign.weights[1][18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold27 (.A(\mydesign.inputs[3][12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mydesign.weights[0][20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mydesign.inputs[3][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mydesign.weights[1][19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mydesign.inputs[3][10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0322_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mydesign.inputs[2][15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0079_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mydesign.inputs[3][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mydesign.inputs[2][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mydesign.weights[2][11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0295_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mydesign.inputs[3][9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0321_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mydesign.weights[2][9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0293_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mydesign.weights[2][19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0012_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mydesign.accum[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0260_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mydesign.inputs[3][15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold48 (.A(\mydesign.inputs[2][10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0015_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mydesign.inputs[2][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold51 (.A(\mydesign.inputs[2][16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mydesign.inputs[3][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mydesign.weights[3][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0113_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mydesign.weights[1][23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mydesign.weights[2][17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0010_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mydesign.weights[2][16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0009_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mydesign.weights[1][17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mydesign.inputs[3][11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0323_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mydesign.inputs[2][17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mydesign.weights[1][16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mydesign.accum[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0188_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mydesign.accum[56] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0220_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mydesign.accum[104] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0124_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mydesign.accum[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0204_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mydesign.weights[2][18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mydesign.weights[1][21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold75 (.A(\mydesign.weights[0][22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mydesign.weights[2][8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0292_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mydesign.inputs[3][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mydesign.weights[0][18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mydesign.weights[1][20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold81 (.A(\mydesign.weights[0][21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mydesign.weights[3][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0114_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mydesign.inputs[2][18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mydesign.inputs[2][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mydesign.weights[3][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0342_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold88 (.A(\mydesign.weights[3][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0115_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mydesign.inputs[3][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0053_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold92 (.A(\mydesign.weights[0][26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mydesign.inputs[3][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0055_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mydesign.weights[0][27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0355_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mydesign.weights[0][25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mydesign.weights[3][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0341_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold100 (.A(\mydesign.inputs[3][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0056_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mydesign.accum[120] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mydesign.weights[0][23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold104 (.A(\mydesign.weights[0][24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0352_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mydesign.weights[3][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0340_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold108 (.A(\mydesign.weights[0][17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mydesign.inputs[0][26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mydesign.accum[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0312_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold112 (.A(\mydesign.weights[3][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0343_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mydesign.weights[2][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mydesign.accum[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0272_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mydesign.inputs[2][19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold118 (.A(\mydesign.weights[1][22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold119 (.A(\mydesign.inputs[0][27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mydesign.accum[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0172_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold122 (.A(\mydesign.weights[2][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mydesign.inputs[3][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0054_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mydesign.cp2[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mydesign.accum[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0236_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mydesign.weights[2][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold129 (.A(\mydesign.weights[0][16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mydesign.accum[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0324_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mydesign.weights[0][19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold133 (.A(\mydesign.weights[2][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mydesign.inputs[0][24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold136 (.A(\mydesign.out[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mydesign.cp2[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mydesign.accum[108] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold139 (.A(\mydesign.accum[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0300_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mydesign.inputs[0][25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold142 (.A(\mydesign.weights[1][14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mydesign.inputs[1][12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mydesign.weights[1][15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold145 (.A(\mydesign.weights[1][13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mydesign.inputs[0][12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold147 (.A(\mydesign.inputs[0][17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold148 (.A(\mydesign.weights[0][12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold149 (.A(\mydesign.inputs[0][21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold150 (.A(\mydesign.inputs[1][13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mydesign.weights[1][10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold152 (.A(\mydesign.weights[1][12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mydesign.inputs[0][14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold154 (.A(\mydesign.accum[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold155 (.A(\mydesign.weights[1][9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold156 (.A(\mydesign.inputs[1][15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold157 (.A(\mydesign.inputs[1][18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold158 (.A(\mydesign.weights[1][11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold159 (.A(\mydesign.inputs[1][19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold160 (.A(\mydesign.inputs[1][21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold161 (.A(\mydesign.inputs[0][16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold162 (.A(\mydesign.weights[0][15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold163 (.A(\mydesign.inputs[1][17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold164 (.A(\mydesign.inputs[0][20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold165 (.A(\mydesign.weights[0][14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mydesign.inputs[0][22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold167 (.A(\mydesign.inputs[0][13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold168 (.A(\mydesign.inputs[0][15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold169 (.A(\mydesign.inputs[0][18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold170 (.A(\mydesign.pe_weights[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0235_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold172 (.A(\mydesign.inputs[1][10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mydesign.inputs[0][23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold174 (.A(\mydesign.inputs[1][22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold175 (.A(\mydesign.inputs[1][8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold176 (.A(\mydesign.inputs[1][20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold177 (.A(\mydesign.inputs[1][16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold178 (.A(\mydesign.inputs[1][14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold179 (.A(\mydesign.inputs[1][23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold180 (.A(\mydesign.inputs[1][9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold181 (.A(\mydesign.inputs[1][11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold182 (.A(\mydesign.inputs[0][19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold183 (.A(\mydesign.weights[1][8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold184 (.A(\mydesign.weights[0][13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold185 (.A(\mydesign.accum[91] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold186 (.A(\mydesign.weights[2][12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold187 (.A(\mydesign.accum[94] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold188 (.A(\mydesign.weights[2][13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold189 (.A(\mydesign.pe_weights[60] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0084_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold191 (.A(\mydesign.weights[2][14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold192 (.A(\mydesign.pe_weights[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0217_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold194 (.A(\mydesign.pe_weights[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0234_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold196 (.A(\mydesign.pe_weights[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold197 (.A(\mydesign.pe_weights[35] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0271_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold199 (.A(\mydesign.accum[57] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0221_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold201 (.A(\mydesign.weights[3][11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold202 (.A(_1776_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0251_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold204 (.A(\mydesign.weights[3][13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold205 (.A(_2507_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0365_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold207 (.A(\mydesign.accum[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold208 (.A(\mydesign.accum[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold209 (.A(\mydesign.pe_weights[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0269_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold211 (.A(\mydesign.pe_weights[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0258_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold213 (.A(\mydesign.pe_inputs[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0310_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold215 (.A(\mydesign.out[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold216 (.A(\mydesign.accum[111] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold217 (.A(\mydesign.pe_inputs[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold218 (.A(\mydesign.accum[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold219 (.A(\mydesign.pe_weights[62] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0154_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold221 (.A(\mydesign.accum[61] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold222 (.A(\mydesign.accum[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold223 (.A(\mydesign.load_counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold224 (.A(\mydesign.accum[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold225 (.A(\mydesign.weights[3][8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold226 (.A(_1770_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0248_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold228 (.A(\mydesign.accum[98] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0142_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold230 (.A(\mydesign.pe_inputs[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0253_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold232 (.A(\mydesign.accum[113] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0105_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold234 (.A(\mydesign.weights[3][10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold235 (.A(_1774_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0250_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold237 (.A(\mydesign.pe_weights[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0233_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold239 (.A(\mydesign.weights[3][9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold240 (.A(_1772_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0249_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold242 (.A(\mydesign.accum[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold243 (.A(\mydesign.pe_weights[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0257_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold245 (.A(\mydesign.accum[35] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold246 (.A(\mydesign.accum[87] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold247 (.A(\mydesign.accum[60] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold248 (.A(\mydesign.compute_en ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold249 (.A(\mydesign.accum[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold250 (.A(\mydesign.weights[3][15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold251 (.A(_2509_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0367_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold253 (.A(\mydesign.pe_weights[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold254 (.A(\mydesign.accum[66] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0206_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold256 (.A(\mydesign.accum[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0189_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold258 (.A(\mydesign.accum[114] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0106_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold260 (.A(\mydesign.pe_inputs[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold261 (.A(\mydesign.pe_weights[61] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold262 (.A(\mydesign.pe_weights[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold263 (.A(\mydesign.accum[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0190_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold265 (.A(\mydesign.accum[62] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold266 (.A(\mydesign.weights[2][15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold267 (.A(\mydesign.accum[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold268 (.A(\mydesign.pe_inputs[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0231_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold270 (.A(\mydesign.accum[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold271 (.A(\mydesign.accum[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold272 (.A(\mydesign.pe_weights[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold273 (.A(\mydesign.accum[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0237_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold275 (.A(\mydesign.accum[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold276 (.A(\mydesign.accum[86] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold277 (.A(\mydesign.accum[89] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0157_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold279 (.A(\mydesign.accum[118] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold280 (.A(\mydesign.pe_inputs[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold281 (.A(\mydesign.accum[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0238_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold283 (.A(\mydesign.accum[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold284 (.A(\mydesign.pe_weights[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0268_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold286 (.A(\mydesign.accum[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold287 (.A(\mydesign.accum[67] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold288 (.A(\mydesign.accum[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0205_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold290 (.A(\mydesign.accum[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold291 (.A(\mydesign.pe_weights[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold292 (.A(\mydesign.accum[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold293 (.A(\mydesign.accum[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold294 (.A(\mydesign.accum[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0274_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold296 (.A(\mydesign.accum[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold297 (.A(\mydesign.accum[105] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0125_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold299 (.A(\mydesign.accum[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold300 (.A(\mydesign.accum[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0273_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold302 (.A(\mydesign.accum[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0262_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold304 (.A(\mydesign.accum[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0286_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold306 (.A(\mydesign.pe_weights[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold307 (.A(\mydesign.accum[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold308 (.A(\mydesign.pe_weights[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold309 (.A(\mydesign.accum[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0313_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold311 (.A(\mydesign.weights[3][14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold312 (.A(_2508_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0366_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold314 (.A(\mydesign.accum[84] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold315 (.A(\mydesign.pe_inputs[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0309_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold317 (.A(\mydesign.accum[115] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold318 (.A(\mydesign.accum[121] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold319 (.A(\mydesign.pe_weights[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold320 (.A(\mydesign.pe_inputs[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold321 (.A(\mydesign.accum[103] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold322 (.A(\mydesign.accum[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold323 (.A(\mydesign.accum[109] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold324 (.A(\mydesign.pe_weights[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold325 (.A(\mydesign.accum[102] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold326 (.A(\mydesign.accum[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold327 (.A(\mydesign.pe_inputs[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0311_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold329 (.A(\mydesign.accum[95] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold330 (.A(\mydesign.accum[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0261_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold332 (.A(\mydesign.accum[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold333 (.A(\mydesign.pe_weights[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0218_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold335 (.A(\mydesign.accum[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0285_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold337 (.A(\mydesign.pe_inputs[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0167_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold339 (.A(\mydesign.accum[122] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold340 (.A(\mydesign.accum[58] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold341 (.A(\mydesign.accum[117] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold342 (.A(\mydesign.accum[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0174_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold344 (.A(\mydesign.accum[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold345 (.A(\mydesign.accum[90] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0158_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold347 (.A(\mydesign.pe_inputs[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold348 (.A(\mydesign.accum[99] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold349 (.A(\mydesign.accum[101] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold350 (.A(\mydesign.accum[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold351 (.A(\mydesign.accum[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold352 (.A(\mydesign.pe_weights[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold353 (.A(\mydesign.accum[116] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold354 (.A(\mydesign.accum[119] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold355 (.A(\mydesign.pe_inputs[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0255_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold357 (.A(\mydesign.pe_inputs[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold358 (.A(\mydesign.accum[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold359 (.A(\mydesign.accum[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold360 (.A(\mydesign.accum[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold361 (.A(\mydesign.accum[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold362 (.A(\mydesign.pe_inputs[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0182_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold364 (.A(\mydesign.accum[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0173_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold366 (.A(\mydesign.weights[3][12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold367 (.A(_2506_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0364_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold369 (.A(\mydesign.pe_weights[58] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold370 (.A(\mydesign.pe_weights[57] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold371 (.A(\mydesign.accum[59] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold372 (.A(\mydesign.accum[112] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold373 (.A(\mydesign.accum[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold374 (.A(\mydesign.pe_inputs[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0183_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold376 (.A(\mydesign.pe_weights[56] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold377 (.A(\mydesign.pe_weights[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold378 (.A(\mydesign.accum[92] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold379 (.A(\mydesign.accum[110] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold380 (.A(\mydesign.accum[93] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold381 (.A(\mydesign.pe_inputs[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0299_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold383 (.A(\mydesign.accum[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold384 (.A(\mydesign.accum[88] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold385 (.A(\mydesign.accum[127] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold386 (.A(\mydesign.accum[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold387 (.A(\mydesign.accum[100] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold388 (.A(\mydesign.accum[97] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0141_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold390 (.A(\mydesign.accum[107] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold391 (.A(\mydesign.accum[106] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0126_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold393 (.A(\mydesign.accum[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold394 (.A(\mydesign.pe_weights[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0232_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold396 (.A(\mydesign.pe_inputs[57] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0097_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold398 (.A(\mydesign.pe_weights[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold399 (.A(\mydesign.accum[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold400 (.A(\mydesign.accum[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold401 (.A(\mydesign.accum[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0302_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold403 (.A(\mydesign.pe_inputs[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0228_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold405 (.A(\mydesign.pe_inputs[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold406 (.A(\mydesign.pe_weights[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0259_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold408 (.A(\mydesign.pe_inputs[58] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0098_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold410 (.A(\mydesign.accum[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0301_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold412 (.A(\mydesign.pe_inputs[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0230_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold414 (.A(\mydesign.pe_weights[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0200_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold416 (.A(\mydesign.accum[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold417 (.A(\mydesign.pe_inputs[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold418 (.A(\mydesign.pe_inputs[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold419 (.A(\mydesign.accum[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0314_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold421 (.A(\mydesign.accum[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold422 (.A(_0326_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold423 (.A(\mydesign.accum[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold424 (.A(\mydesign.pe_weights[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold425 (.A(\mydesign.load_counter[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold426 (.A(\mydesign.accum[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold427 (.A(\mydesign.pe_inputs[59] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0119_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold429 (.A(\mydesign.accum[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold430 (.A(\mydesign.accum[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold431 (.A(\mydesign.pe_inputs[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0164_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold433 (.A(\mydesign.accum[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold434 (.A(\mydesign.accum[96] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0937_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold436 (.A(\mydesign.accum[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold437 (.A(_0319_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold438 (.A(\mydesign.accum[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0325_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold440 (.A(\mydesign.pe_inputs[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold441 (.A(\mydesign.accum[125] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold442 (.A(\mydesign.accum[123] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold443 (.A(\mydesign.accum[126] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold444 (.A(\mydesign.accum[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold445 (.A(\mydesign.load_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold446 (.A(\mydesign.pe_inputs[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0308_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold448 (.A(\mydesign.pe_weights[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold449 (.A(\mydesign.accum[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold450 (.A(net9),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold451 (.A(_0069_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold452 (.A(\mydesign.pe_inputs[61] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold453 (.A(net14),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold454 (.A(\mydesign.pe_inputs[56] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold455 (.A(_0096_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold456 (.A(net12),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold457 (.A(\mydesign.pe_inputs[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold458 (.A(\mydesign.pe_weights[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold459 (.A(net11),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold460 (.A(\mydesign.accum[124] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold461 (.A(net13),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold462 (.A(net8),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold463 (.A(\mydesign.pe_inputs[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold464 (.A(\mydesign.cp[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold465 (.A(net15),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0075_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold467 (.A(\mydesign.pe_inputs[62] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold468 (.A(net10),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold469 (.A(\mydesign.cp[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold470 (.A(\mydesign.accum[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold471 (.A(\mydesign.pe_inputs[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold472 (.A(\mydesign.pe_weights[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold473 (.A(\mydesign.pe_weights[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold474 (.A(\mydesign.load_counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold475 (.A(\mydesign.pe_inputs[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold476 (.A(\mydesign.pe_inputs[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold477 (.A(\mydesign.pe_weights[59] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold478 (.A(\mydesign.pe_inputs[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold479 (.A(\mydesign.pe_inputs[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0296_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold481 (.A(\mydesign.pe_inputs[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold482 (.A(\mydesign.pe_weights[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold483 (.A(\mydesign.pe_inputs[60] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold484 (.A(\mydesign.out[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold485 (.A(_0339_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold486 (.A(\mydesign.out[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold487 (.A(\mydesign.load_counter[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold488 (.A(\mydesign.pe_inputs[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold489 (.A(\mydesign.load_counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold490 (.A(_2639_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold491 (.A(\mydesign.load_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold492 (.A(\mydesign.pe_inputs[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1111));
 sg13g2_decap_4 FILLER_0_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net399;
 assign uio_oe[1] = net400;
 assign uio_oe[2] = net401;
 assign uio_oe[3] = net402;
 assign uio_oe[4] = net403;
 assign uio_oe[5] = net404;
 assign uio_oe[6] = net405;
 assign uio_oe[7] = net406;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
endmodule
